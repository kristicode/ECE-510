*** SPICE deck for cell testJTLplain{sch} from library aNewTestLibrary
*** Created on Sat Jan 09, 2021 14:13:09
*** Last revised on Mon Aug 26, 2024 11:38:12
*** Written on Mon Aug 26, 2024 11:55:08 by Electric VLSI Design System, version 9.08e
*** Layout tech: josephson, foundry NONE
*** UC SPICE *** , MIN_RESIST 0.0, MIN_CAPAC 0.0FF
* Model cards copied from file: /Users/ivans/years/2020-2024/2024/2024-ivan/electric-2024/theBest1aug24/aTests/testJTLplain.txt
*** These are the print statement for testJTLplain
*** ies 26 August 2024
*** josim -o Aoutput.csv testJTLplain.cir 



.tran 0.1p 20p 0 0.1p


.print DEVV BJi|xJ28
.print DEVV BJi|xJ37
.print DEVV BJi|xJ64
.print DEVV BJi|xJ73




* End of Model cards copied from file: /Users/ivans/years/2020-2024/2024/2024-ivan/electric-2024/theBest1jul24/aTests/testJTL.txt
.model jmitll jj(rtype=1, vg=.002V, cap=0.07pF, r0=160, rN=16, icrit=0.0001A)


.SUBCKT junctionsBypassGround__gbj1p0 D 
BJi D gnd jmitll area=1.25
RRi D gnd 5.36
.ENDS junctionsBypassGround__gbj1p0


*** SUBCIRCUIT inductors__fixedInd1p5 FROM CELL inductors:fixedInd3p0{sch}
.SUBCKT inductors__fixedInd1p5 A B
LLi A B 7.891E-12
.ENDS inductors__fixedInd1p5


*** SUBCIRCUIT conductors__anyBias-Lk_0 FROM CELL conductors:anyBias{sch}
.SUBCKT conductors__anyBias-Lk_0  D
RR1 NN D 29.42
VrampSppl@0 NN gnd pwl (0 0 1p 0.0026V)
.ENDS conductors__anyBias-Lk_0_707



****.SUBCKT conductors__anyBias-Lk_0 D
****RR1 NN D 8
****VrampSppl@0 NN gnd pwl (0 0 1p 3.86V)
***.ENDS conductors__anyBias-Lk_0

*** SUBCIRCUIT junctions__jb2p0 FROM CELL junctions:jb2p0{sch}
.SUBCKT junctions__jb2p0 D S
BJi S D jmitll area=2.5
RRi S D 2.68
.ENDS junctions__jb2p0

*** SUBCIRCUIT junctions__jb200p0 FROM CELL junctions:jb200p0{sch}
.SUBCKT junctions__jb200p0 D S
BJi S D jmitll area=250.0
RRi S D 0.0268
.ENDS junctions__jb200p0

*** SUBCIRCUIT conductors__anyBias-Lk_1_414 FROM CELL conductors:anyBias{sch}
.SUBCKT conductors__anyBias-Lk_1_414 D
RR1 NN D 14.71
VrampSppl@0 NN gnd pwl (0 0 1p 0.0026V)
.ENDS conductors__anyBias-Lk_1_414

*** SUBCIRCUIT conductors__bias1p4 FROM CELL conductors:bias1p4{sch}
.SUBCKT conductors__bias1p4 D
Xnormaliz@0 D conductors__anyBias-Lk_1_414
.ENDS conductors__bias1p4

*** SUBCIRCUIT conductors__anyBias-Lk_141_4 FROM CELL conductors:anyBias{sch}
.SUBCKT conductors__anyBias-Lk_141_4 D
RR1 NN D 0.147
VrampSppl@0 NN gnd pwl (0 0 1p 0.0026V)
.ENDS conductors__anyBias-Lk_141_4

*** SUBCIRCUIT conductors__bias1p4x100 FROM CELL conductors:bias1p4x100{sch}
.SUBCKT conductors__bias1p4x100 D
Xnormaliz@0 D conductors__anyBias-Lk_141_4
.ENDS conductors__bias1p4x100

*** SUBCIRCUIT newJTL__phaseReference FROM CELL newJTL:phaseReference{sch}
.SUBCKT newJTL__phaseReference B1 B2 gnd
XJ1 gnd B1 junctions__jb2p0
XJ2 gnd B2 junctions__jb200p0
LM1 net@4 B1 10e-16
LM2 net@3 B2 10e-16
Xbias1p4@0 net@4 conductors__bias1p4
Xbias1p4x@0 net@3 conductors__bias1p4x100
.ENDS newJTL__phaseReference



**cart_pole_input**
.SUBCKT conductors__anyBias-Lk_0_701 bottom out
VrampSppl@0 bottom out pwl(8000p 1mV 8001p 0mV 13000p 1mV 13001p 0mV 22000p 1mV 22001p 0mV 44000p 1mV 44001p 0mV 52000p 1mV 52001p 0mV 55000p 1mV 55001p 0mV 83000p 1mV 83001p 0mV 87000p 1mV 87001p 0mV 91000p 1mV 91001p 0mV 115000p 1mV 115001p 0mV 121000p 1mV 121001p 0mV 137000p 1mV 137001p 0mV 140000p 1mV 140001p 0mV 141000p 1mV 141001p 0mV 188000p 1mV 188001p 0mV 204000p 1mV 204001p 0mV 219000p 1mV 219001p 0mV 226000p 1mV 226001p 0mV 229000p 1mV 229001p 0mV 233000p 1mV 233001p 0mV 249000p 1mV 249001p 0mV 254000p 1mV 254001p 0mV 259000p 1mV 259001p 0mV 268000p 1mV 268001p 0mV 281000p 1mV 281001p 0mV 301000p 1mV 301001p 0mV 302000p 1mV 302001p 0mV 313000p 1mV 313001p 0mV 339000p 1mV 339001p 0mV 346000p 1mV 346001p 0mV 381000p 1mV 381001p 0mV 396000p 1mV 396001p 0mV 410000p 1mV 410001p 0mV 436000p 1mV 436001p 0mV 452000p 1mV 452001p 0mV 456000p 1mV 456001p 0mV 476000p 1mV 476001p 0mV 484000p 1mV 484001p 0mV 486000p 1mV 486001p 0mV 495000p 1mV 495001p 0mV 496000p 1mV 496001p 0mV 513000p 1mV 513001p 0mV 542000p 1mV 542001p 0mV 543000p 1mV 543001p 0mV 625000p 1mV 625001p 0mV 650000p 1mV 650001p 0mV 712000p 1mV 712001p 0mV 734000p 1mV 734001p 0mV 767000p 1mV 767001p 0mV 771000p 1mV 771001p 0mV 777000p 1mV 777001p 0mV 780000p 1mV 780001p 0mV 804000p 1mV 804001p 0mV 813000p 1mV 813001p 0mV 829000p 1mV 829001p 0mV 830000p 1mV 830001p 0mV 836000p 1mV 836001p 0mV 838000p 1mV 838001p 0mV 839000p 1mV 839001p 0mV 862000p 1mV 862001p 0mV 890000p 1mV 890001p 0mV 894000p 1mV 894001p 0mV 935000p 1mV 935001p 0mV 952000p 1mV 952001p 0mV 954000p 1mV 954001p 0mV 984000p 1mV 984001p 0mV 985000p 1mV 985001p 0mV 1000000p 1mV 1000001p 0mV 1019000p 1mV 1019001p 0mV 1033000p 1mV 1033001p 0mV 1051000p 1mV 1051001p 0mV 1056000p 1mV 1056001p 0mV 1057000p 1mV 1057001p 0mV 1086000p 1mV 1086001p 0mV 1090000p 1mV 1090001p 0mV 1109000p 1mV 1109001p 0mV 1116000p 1mV 1116001p 0mV 1126000p 1mV 1126001p 0mV 1149000p 1mV 1149001p 0mV 1152000p 1mV 1152001p 0mV 1276000p 1mV 1276001p 0mV 1287000p 1mV 1287001p 0mV 1311000p 1mV 1311001p 0mV 1315000p 1mV 1315001p 0mV 1323000p 1mV 1323001p 0mV 1328000p 1mV 1328001p 0mV 1354000p 1mV 1354001p 0mV 1359000p 1mV 1359001p 0mV 1375000p 1mV 1375001p 0mV 1382000p 1mV 1382001p 0mV 1397000p 1mV 1397001p 0mV 1419000p 1mV 1419001p 0mV 1452000p 1mV 1452001p 0mV 1455000p 1mV 1455001p 0mV 1490000p 1mV 1490001p 0mV 1522000p 1mV 1522001p 0mV 1561000p 1mV 1561001p 0mV 1571000p 1mV 1571001p 0mV 1578000p 1mV 1578001p 0mV 1583000p 1mV 1583001p 0mV 1598000p 1mV 1598001p 0mV 1609000p 1mV 1609001p 0mV 1633000p 1mV 1633001p 0mV 1658000p 1mV 1658001p 0mV 1671000p 1mV 1671001p 0mV 1740000p 1mV 1740001p 0mV 1754000p 1mV 1754001p 0mV 1763000p 1mV 1763001p 0mV 1771000p 1mV 1771001p 0mV 1787000p 1mV 1787001p 0mV 1797000p 1mV 1797001p 0mV 1808000p 1mV 1808001p 0mV 1810000p 1mV 1810001p 0mV 1838000p 1mV 1838001p 0mV 1841000p 1mV 1841001p 0mV 1850000p 1mV 1850001p 0mV 1854000p 1mV 1854001p 0mV 1873000p 1mV 1873001p 0mV 1884000p 1mV 1884001p 0mV 1887000p 1mV 1887001p 0mV 1897000p 1mV 1897001p 0mV 1901000p 1mV 1901001p 0mV 1903000p 1mV 1903001p 0mV 1928000p 1mV 1928001p 0mV 1933000p 1mV 1933001p 0mV 1961000p 1mV 1961001p 0mV 1978000p 1mV 1978001p 0mV 1980000p 1mV 1980001p 0mV 2003000p 1mV 2003001p 0mV 2020000p 1mV 2020001p 0mV 2028000p 1mV 2028001p 0mV 2030000p 1mV 2030001p 0mV 2039000p 1mV 2039001p 0mV 2048000p 1mV 2048001p 0mV 2056000p 1mV 2056001p 0mV 2081000p 1mV 2081001p 0mV 2090000p 1mV 2090001p 0mV 2115000p 1mV 2115001p 0mV 2124000p 1mV 2124001p 0mV 2126000p 1mV 2126001p 0mV 2157000p 1mV 2157001p 0mV 2164000p 1mV 2164001p 0mV 2173000p 1mV 2173001p 0mV 2174000p 1mV 2174001p 0mV 2200000p 1mV 2200001p 0mV 2209000p 1mV 2209001p 0mV 2220000p 1mV 2220001p 0mV 2228000p 1mV 2228001p 0mV 2231000p 1mV 2231001p 0mV 2233000p 1mV 2233001p 0mV 2239000p 1mV 2239001p 0mV 2333000p 1mV 2333001p 0mV 2335000p 1mV 2335001p 0mV 2338000p 1mV 2338001p 0mV 2355000p 1mV 2355001p 0mV 2387000p 1mV 2387001p 0mV 2390000p 1mV 2390001p 0mV 2418000p 1mV 2418001p 0mV 2421000p 1mV 2421001p 0mV 2427000p 1mV 2427001p 0mV 2501000p 1mV 2501001p 0mV 2548000p 1mV 2548001p 0mV 2558000p 1mV 2558001p 0mV 2584000p 1mV 2584001p 0mV 2589000p 1mV 2589001p 0mV 2641000p 1mV 2641001p 0mV 2665000p 1mV 2665001p 0mV 2682000p 1mV 2682001p 0mV 2712000p 1mV 2712001p 0mV 2740000p 1mV 2740001p 0mV 2766000p 1mV 2766001p 0mV 2775000p 1mV 2775001p 0mV 2818000p 1mV 2818001p 0mV 2842000p 1mV 2842001p 0mV 2858000p 1mV 2858001p 0mV 2888000p 1mV 2888001p 0mV 2903000p 1mV 2903001p 0mV 2913000p 1mV 2913001p 0mV 2983000p 1mV 2983001p 0mV 2989000p 1mV 2989001p 0mV 3035000p 1mV 3035001p 0mV 3054000p 1mV 3054001p 0mV 3113000p 1mV 3113001p 0mV 3136000p 1mV 3136001p 0mV 3163000p 1mV 3163001p 0mV 3166000p 1mV 3166001p 0mV 3174000p 1mV 3174001p 0mV 3175000p 1mV 3175001p 0mV 3186000p 1mV 3186001p 0mV 3207000p 1mV 3207001p 0mV 3238000p 1mV 3238001p 0mV 3256000p 1mV 3256001p 0mV 3258000p 1mV 3258001p 0mV 3264000p 1mV 3264001p 0mV 3276000p 1mV 3276001p 0mV 3280000p 1mV 3280001p 0mV 3292000p 1mV 3292001p 0mV 3308000p 1mV 3308001p 0mV 3392000p 1mV 3392001p 0mV 3410000p 1mV 3410001p 0mV 3419000p 1mV 3419001p 0mV 3445000p 1mV 3445001p 0mV 3446000p 1mV 3446001p 0mV 3458000p 1mV 3458001p 0mV 3464000p 1mV 3464001p 0mV 3479000p 1mV 3479001p 0mV 3515000p 1mV 3515001p 0mV 3520000p 1mV 3520001p 0mV 3522000p 1mV 3522001p 0mV 3525000p 1mV 3525001p 0mV 3542000p 1mV 3542001p 0mV 3565000p 1mV 3565001p 0mV 3585000p 1mV 3585001p 0mV 3611000p 1mV 3611001p 0mV 3640000p 1mV 3640001p 0mV 3666000p 1mV 3666001p 0mV 3681000p 1mV 3681001p 0mV 3682000p 1mV 3682001p 0mV 3706000p 1mV 3706001p 0mV 3739000p 1mV 3739001p 0mV 3742000p 1mV 3742001p 0mV 3744000p 1mV 3744001p 0mV 3755000p 1mV 3755001p 0mV 3766000p 1mV 3766001p 0mV 3775000p 1mV 3775001p 0mV 3778000p 1mV 3778001p 0mV 3861000p 1mV 3861001p 0mV 3908000p 1mV 3908001p 0mV 3917000p 1mV 3917001p 0mV 3921000p 1mV 3921001p 0mV 3929000p 1mV 3929001p 0mV 3936000p 1mV 3936001p 0mV 3944000p 1mV 3944001p 0mV 3953000p 1mV 3953001p 0mV 3956000p 1mV 3956001p 0mV 3965000p 1mV 3965001p 0mV 3994000p 1mV 3994001p 0mV 4021000p 1mV 4021001p 0mV 4026000p 1mV 4026001p 0mV 4027000p 1mV 4027001p 0mV 4031000p 1mV 4031001p 0mV 4046000p 1mV 4046001p 0mV 4056000p 1mV 4056001p 0mV 4063000p 1mV 4063001p 0mV 4095000p 1mV 4095001p 0mV 4098000p 1mV 4098001p 0mV 4106000p 1mV 4106001p 0mV 4133000p 1mV 4133001p 0mV 4155000p 1mV 4155001p 0mV 4158000p 1mV 4158001p 0mV 4169000p 1mV 4169001p 0mV 4179000p 1mV 4179001p 0mV 4236000p 1mV 4236001p 0mV 4248000p 1mV 4248001p 0mV 4253000p 1mV 4253001p 0mV 4268000p 1mV 4268001p 0mV 4271000p 1mV 4271001p 0mV 4276000p 1mV 4276001p 0mV 4282000p 1mV 4282001p 0mV 4336000p 1mV 4336001p 0mV 4360000p 1mV 4360001p 0mV 4363000p 1mV 4363001p 0mV 4367000p 1mV 4367001p 0mV 4368000p 1mV 4368001p 0mV 4369000p 1mV 4369001p 0mV 4374000p 1mV 4374001p 0mV 4384000p 1mV 4384001p 0mV 4418000p 1mV 4418001p 0mV 4429000p 1mV 4429001p 0mV 4457000p 1mV 4457001p 0mV 4462000p 1mV 4462001p 0mV 4463000p 1mV 4463001p 0mV 4470000p 1mV 4470001p 0mV 4483000p 1mV 4483001p 0mV 4485000p 1mV 4485001p 0mV 4497000p 1mV 4497001p 0mV 4516000p 1mV 4516001p 0mV 4520000p 1mV 4520001p 0mV 4523000p 1mV 4523001p 0mV 4532000p 1mV 4532001p 0mV 4550000p 1mV 4550001p 0mV 4552000p 1mV 4552001p 0mV 4557000p 1mV 4557001p 0mV 4563000p 1mV 4563001p 0mV 4578000p 1mV 4578001p 0mV 4586000p 1mV 4586001p 0mV 4606000p 1mV 4606001p 0mV 4614000p 1mV 4614001p 0mV 4619000p 1mV 4619001p 0mV 4670000p 1mV 4670001p 0mV 4716000p 1mV 4716001p 0mV 4718000p 1mV 4718001p 0mV 4741000p 1mV 4741001p 0mV 4765000p 1mV 4765001p 0mV 4768000p 1mV 4768001p 0mV 4770000p 1mV 4770001p 0mV 4772000p 1mV 4772001p 0mV 4780000p 1mV 4780001p 0mV 4828000p 1mV 4828001p 0mV 4835000p 1mV 4835001p 0mV 4852000p 1mV 4852001p 0mV 4859000p 1mV 4859001p 0mV 4872000p 1mV 4872001p 0mV 4878000p 1mV 4878001p 0mV 4902000p 1mV 4902001p 0mV 4903000p 1mV 4903001p 0mV 4912000p 1mV 4912001p 0mV 4914000p 1mV 4914001p 0mV 4915000p 1mV 4915001p 0mV 4931000p 1mV 4931001p 0mV 4935000p 1mV 4935001p 0mV 4939000p 1mV 4939001p 0mV 4953000p 1mV 4953001p 0mV 4978000p 1mV 4978001p 0mV 4992000p 1mV 4992001p 0mV 5019000p 1mV 5019001p 0mV 5028000p 1mV 5028001p 0mV 5036000p 1mV 5036001p 0mV 5046000p 1mV 5046001p 0mV 5068000p 1mV 5068001p 0mV 5078000p 1mV 5078001p 0mV 5104000p 1mV 5104001p 0mV 5110000p 1mV 5110001p 0mV 5112000p 1mV 5112001p 0mV 5122000p 1mV 5122001p 0mV 5126000p 1mV 5126001p 0mV 5138000p 1mV 5138001p 0mV 5146000p 1mV 5146001p 0mV 5158000p 1mV 5158001p 0mV 5161000p 1mV 5161001p 0mV 5166000p 1mV 5166001p 0mV 5180000p 1mV 5180001p 0mV 5195000p 1mV 5195001p 0mV 5240000p 1mV 5240001p 0mV 5242000p 1mV 5242001p 0mV 5259000p 1mV 5259001p 0mV 5271000p 1mV 5271001p 0mV 5277000p 1mV 5277001p 0mV 5293000p 1mV 5293001p 0mV 5308000p 1mV 5308001p 0mV 5310000p 1mV 5310001p 0mV 5317000p 1mV 5317001p 0mV 5328000p 1mV 5328001p 0mV 5339000p 1mV 5339001p 0mV 5351000p 1mV 5351001p 0mV 5352000p 1mV 5352001p 0mV 5367000p 1mV 5367001p 0mV 5369000p 1mV 5369001p 0mV 5383000p 1mV 5383001p 0mV 5396000p 1mV 5396001p 0mV 5412000p 1mV 5412001p 0mV 5414000p 1mV 5414001p 0mV 5455000p 1mV 5455001p 0mV 5456000p 1mV 5456001p 0mV 5511000p 1mV 5511001p 0mV 5519000p 1mV 5519001p 0mV 5535000p 1mV 5535001p 0mV 5573000p 1mV 5573001p 0mV 5598000p 1mV 5598001p 0mV 5605000p 1mV 5605001p 0mV 5644000p 1mV 5644001p 0mV 5661000p 1mV 5661001p 0mV 5752000p 1mV 5752001p 0mV 5767000p 1mV 5767001p 0mV 5799000p 1mV 5799001p 0mV 5825000p 1mV 5825001p 0mV 5847000p 1mV 5847001p 0mV 5850000p 1mV 5850001p 0mV 5857000p 1mV 5857001p 0mV 5864000p 1mV 5864001p 0mV 5867000p 1mV 5867001p 0mV 5881000p 1mV 5881001p 0mV 5923000p 1mV 5923001p 0mV 5927000p 1mV 5927001p 0mV 5928000p 1mV 5928001p 0mV 5985000p 1mV 5985001p 0mV 6000000p 1mV 6000001p 0mV 6037000p 1mV 6037001p 0mV 6039000p 1mV 6039001p 0mV 6075000p 1mV 6075001p 0mV 6092000p 1mV 6092001p 0mV 6096000p 1mV 6096001p 0mV 6116000p 1mV 6116001p 0mV 6128000p 1mV 6128001p 0mV 6162000p 1mV 6162001p 0mV 6168000p 1mV 6168001p 0mV 6192000p 1mV 6192001p 0mV 6237000p 1mV 6237001p 0mV 6247000p 1mV 6247001p 0mV 6258000p 1mV 6258001p 0mV 6286000p 1mV 6286001p 0mV 6293000p 1mV 6293001p 0mV 6300000p 1mV 6300001p 0mV 6362000p 1mV 6362001p 0mV 6408000p 1mV 6408001p 0mV 6492000p 1mV 6492001p 0mV 6520000p 1mV 6520001p 0mV 6539000p 1mV 6539001p 0mV 6551000p 1mV 6551001p 0mV 6565000p 1mV 6565001p 0mV 6574000p 1mV 6574001p 0mV 6608000p 1mV 6608001p 0mV 6620000p 1mV 6620001p 0mV 6631000p 1mV 6631001p 0mV 6663000p 1mV 6663001p 0mV 6674000p 1mV 6674001p 0mV 6677000p 1mV 6677001p 0mV 6802000p 1mV 6802001p 0mV 6803000p 1mV 6803001p 0mV 6821000p 1mV 6821001p 0mV 6829000p 1mV 6829001p 0mV 6863000p 1mV 6863001p 0mV 7032000p 1mV 7032001p 0mV 7050000p 1mV 7050001p 0mV 7234000p 1mV 7234001p 0mV 7283000p 1mV 7283001p 0mV 7431000p 1mV 7431001p 0mV 7508000p 1mV 7508001p 0mV 7616000p 1mV 7616001p 0mV 7643000p 1mV 7643001p 0mV 7656000p 1mV 7656001p 0mV 7664000p 1mV 7664001p 0mV 7914000p 1mV 7914001p 0mV 7984000p 1mV 7984001p 0mV 8048000p 1mV 8048001p 0mV 8051000p 1mV 8051001p 0mV 8220000p 1mV 8220001p 0mV 8258000p 1mV 8258001p 0mV 8277000p 1mV 8277001p 0mV 8311000p 1mV 8311001p 0mV 8329000p 1mV 8329001p 0mV 8379000p 1mV 8379001p 0mV 8385000p 1mV 8385001p 0mV 8394000p 1mV 8394001p 0mV 8447000p 1mV 8447001p 0mV 8461000p 1mV 8461001p 0mV 8540000p 1mV 8540001p 0mV 8600000p 1mV 8600001p 0mV 8663000p 1mV 8663001p 0mV 8665000p 1mV 8665001p 0mV 8669000p 1mV 8669001p 0mV 8720000p 1mV 8720001p 0mV 8800000p 1mV 8800001p 0mV 8816000p 1mV 8816001p 0mV 8833000p 1mV 8833001p 0mV 8849000p 1mV 8849001p 0mV 8866000p 1mV 8866001p 0mV 8959000p 1mV 8959001p 0mV 9011000p 1mV 9011001p 0mV 9013000p 1mV 9013001p 0mV 9073000p 1mV 9073001p 0mV 9077000p 1mV 9077001p 0mV 9146000p 1mV 9146001p 0mV 9165000p 1mV 9165001p 0mV 9204000p 1mV 9204001p 0mV 9208000p 1mV 9208001p 0mV 9298000p 1mV 9298001p 0mV 9434000p 1mV 9434001p 0mV 9459000p 1mV 9459001p 0mV 9700000p 1mV 9700001p 0mV 9731000p 1mV 9731001p 0mV 9732000p 1mV 9732001p 0mV 9791000p 1mV 9791001p 0mV 9794000p 1mV 9794001p 0mV 9805000p 1mV 9805001p 0mV 9854000p 1mV 9854001p 0mV 9897000p 1mV 9897001p 0mV 9899000p 1mV 9899001p 0mV 9903000p 1mV 9903001p 0mV 9934000p 1mV 9934001p 0mV 9942000p 1mV 9942001p 0mV 9949000p 1mV 9949001p 0mV 9987000p 1mV 9987001p 0mV 9998000p 1mV 9998001p 0mV)
.ENDS conductors__anyBias-Lk_0_701


.SUBCKT conductors__anyBias-Lk_0_702 bottom out
VrampSppl@0 bottom out pwl (301000p 1mV 301001p 0mV 302000p 1mV 302001p 0mV 308000p 1mV 308001p 0mV 310000p 1mV 310001p 0mV 311000p 1mV 311001p 0mV 315000p 1mV 315001p 0mV 321000p 1mV 321001p 0mV 337000p 1mV 337001p 0mV 340000p 1mV 340001p 0mV 355000p 1mV 355001p 0mV 362000p 1mV 362001p 0mV 366000p 1mV 366001p 0mV 377000p 1mV 377001p 0mV 378000p 1mV 378001p 0mV 388000p 1mV 388001p 0mV 413000p 1mV 413001p 0mV 424000p 1mV 424001p 0mV 442000p 1mV 442001p 0mV 453000p 1mV 453001p 0mV 456000p 1mV 456001p 0mV 474000p 1mV 474001p 0mV 478000p 1mV 478001p 0mV 487000p 1mV 487001p 0mV 523000p 1mV 523001p 0mV 528000p 1mV 528001p 0mV 553000p 1mV 553001p 0mV 569000p 1mV 569001p 0mV 571000p 1mV 571001p 0mV 602000p 1mV 602001p 0mV 621000p 1mV 621001p 0mV 623000p 1mV 623001p 0mV 624000p 1mV 624001p 0mV 628000p 1mV 628001p 0mV 633000p 1mV 633001p 0mV 635000p 1mV 635001p 0mV 651000p 1mV 651001p 0mV 656000p 1mV 656001p 0mV 660000p 1mV 660001p 0mV 667000p 1mV 667001p 0mV 675000p 1mV 675001p 0mV 680000p 1mV 680001p 0mV 681000p 1mV 681001p 0mV 682000p 1mV 682001p 0mV 691000p 1mV 691001p 0mV 713000p 1mV 713001p 0mV 718000p 1mV 718001p 0mV 722000p 1mV 722001p 0mV 744000p 1mV 744001p 0mV 746000p 1mV 746001p 0mV 754000p 1mV 754001p 0mV 775000p 1mV 775001p 0mV 780000p 1mV 780001p 0mV 790000p 1mV 790001p 0mV 795000p 1mV 795001p 0mV 798000p 1mV 798001p 0mV 805000p 1mV 805001p 0mV 824000p 1mV 824001p 0mV 826000p 1mV 826001p 0mV 836000p 1mV 836001p 0mV 842000p 1mV 842001p 0mV 848000p 1mV 848001p 0mV 851000p 1mV 851001p 0mV 857000p 1mV 857001p 0mV 861000p 1mV 861001p 0mV 875000p 1mV 875001p 0mV 876000p 1mV 876001p 0mV 879000p 1mV 879001p 0mV 884000p 1mV 884001p 0mV 889000p 1mV 889001p 0mV 896000p 1mV 896001p 0mV 905000p 1mV 905001p 0mV 911000p 1mV 911001p 0mV 915000p 1mV 915001p 0mV 919000p 1mV 919001p 0mV 924000p 1mV 924001p 0mV 928000p 1mV 928001p 0mV 932000p 1mV 932001p 0mV 935000p 1mV 935001p 0mV 979000p 1mV 979001p 0mV 986000p 1mV 986001p 0mV 991000p 1mV 991001p 0mV 1001000p 1mV 1001001p 0mV 1004000p 1mV 1004001p 0mV 1024000p 1mV 1024001p 0mV 1038000p 1mV 1038001p 0mV 1051000p 1mV 1051001p 0mV 1052000p 1mV 1052001p 0mV 1059000p 1mV 1059001p 0mV 1063000p 1mV 1063001p 0mV 1064000p 1mV 1064001p 0mV 1075000p 1mV 1075001p 0mV 1089000p 1mV 1089001p 0mV 1091000p 1mV 1091001p 0mV 1119000p 1mV 1119001p 0mV 1128000p 1mV 1128001p 0mV 1129000p 1mV 1129001p 0mV 1130000p 1mV 1130001p 0mV 1132000p 1mV 1132001p 0mV 1138000p 1mV 1138001p 0mV 1143000p 1mV 1143001p 0mV 1172000p 1mV 1172001p 0mV 1178000p 1mV 1178001p 0mV 1188000p 1mV 1188001p 0mV 1192000p 1mV 1192001p 0mV 1206000p 1mV 1206001p 0mV 1207000p 1mV 1207001p 0mV 1210000p 1mV 1210001p 0mV 1220000p 1mV 1220001p 0mV 1226000p 1mV 1226001p 0mV 1227000p 1mV 1227001p 0mV 1244000p 1mV 1244001p 0mV 1249000p 1mV 1249001p 0mV 1253000p 1mV 1253001p 0mV 1267000p 1mV 1267001p 0mV 1268000p 1mV 1268001p 0mV 1302000p 1mV 1302001p 0mV 1323000p 1mV 1323001p 0mV 1324000p 1mV 1324001p 0mV 1337000p 1mV 1337001p 0mV 1353000p 1mV 1353001p 0mV 1360000p 1mV 1360001p 0mV 1369000p 1mV 1369001p 0mV 1372000p 1mV 1372001p 0mV 1373000p 1mV 1373001p 0mV 1374000p 1mV 1374001p 0mV 1383000p 1mV 1383001p 0mV 1392000p 1mV 1392001p 0mV 1394000p 1mV 1394001p 0mV 1395000p 1mV 1395001p 0mV 1398000p 1mV 1398001p 0mV 1428000p 1mV 1428001p 0mV 1435000p 1mV 1435001p 0mV 1438000p 1mV 1438001p 0mV 1460000p 1mV 1460001p 0mV 1472000p 1mV 1472001p 0mV 1474000p 1mV 1474001p 0mV 1492000p 1mV 1492001p 0mV 1493000p 1mV 1493001p 0mV 1500000p 1mV 1500001p 0mV 1501000p 1mV 1501001p 0mV 1502000p 1mV 1502001p 0mV 1519000p 1mV 1519001p 0mV 1533000p 1mV 1533001p 0mV 1545000p 1mV 1545001p 0mV 1547000p 1mV 1547001p 0mV 1548000p 1mV 1548001p 0mV 1570000p 1mV 1570001p 0mV 1597000p 1mV 1597001p 0mV 1705000p 1mV 1705001p 0mV 1707000p 1mV 1707001p 0mV 1720000p 1mV 1720001p 0mV 1728000p 1mV 1728001p 0mV 1730000p 1mV 1730001p 0mV 1732000p 1mV 1732001p 0mV 1738000p 1mV 1738001p 0mV 1746000p 1mV 1746001p 0mV 1754000p 1mV 1754001p 0mV 1765000p 1mV 1765001p 0mV 1768000p 1mV 1768001p 0mV 1783000p 1mV 1783001p 0mV 1796000p 1mV 1796001p 0mV 1907000p 1mV 1907001p 0mV 1909000p 1mV 1909001p 0mV 1924000p 1mV 1924001p 0mV 1927000p 1mV 1927001p 0mV 1940000p 1mV 1940001p 0mV 1944000p 1mV 1944001p 0mV 1952000p 1mV 1952001p 0mV 1954000p 1mV 1954001p 0mV 1961000p 1mV 1961001p 0mV 1968000p 1mV 1968001p 0mV 1973000p 1mV 1973001p 0mV 1979000p 1mV 1979001p 0mV 1994000p 1mV 1994001p 0mV 2103000p 1mV 2103001p 0mV 2106000p 1mV 2106001p 0mV 2116000p 1mV 2116001p 0mV 2125000p 1mV 2125001p 0mV 2130000p 1mV 2130001p 0mV 2152000p 1mV 2152001p 0mV 2153000p 1mV 2153001p 0mV 2159000p 1mV 2159001p 0mV 2160000p 1mV 2160001p 0mV 2164000p 1mV 2164001p 0mV 2166000p 1mV 2166001p 0mV 2169000p 1mV 2169001p 0mV 2174000p 1mV 2174001p 0mV 3107000p 1mV 3107001p 0mV 3118000p 1mV 3118001p 0mV 3120000p 1mV 3120001p 0mV 3127000p 1mV 3127001p 0mV 3129000p 1mV 3129001p 0mV 3130000p 1mV 3130001p 0mV 3147000p 1mV 3147001p 0mV 3150000p 1mV 3150001p 0mV 3152000p 1mV 3152001p 0mV 3180000p 1mV 3180001p 0mV 3182000p 1mV 3182001p 0mV 3197000p 1mV 3197001p 0mV 3208000p 1mV 3208001p 0mV 3223000p 1mV 3223001p 0mV 3242000p 1mV 3242001p 0mV 3245000p 1mV 3245001p 0mV 3247000p 1mV 3247001p 0mV 3259000p 1mV 3259001p 0mV 3267000p 1mV 3267001p 0mV 3274000p 1mV 3274001p 0mV 3287000p 1mV 3287001p 0mV 3293000p 1mV 3293001p 0mV 3301000p 1mV 3301001p 0mV 3304000p 1mV 3304001p 0mV 3308000p 1mV 3308001p 0mV 3310000p 1mV 3310001p 0mV 3323000p 1mV 3323001p 0mV 3341000p 1mV 3341001p 0mV 3343000p 1mV 3343001p 0mV 3345000p 1mV 3345001p 0mV 3346000p 1mV 3346001p 0mV 3350000p 1mV 3350001p 0mV 3353000p 1mV 3353001p 0mV 3355000p 1mV 3355001p 0mV 3370000p 1mV 3370001p 0mV 3378000p 1mV 3378001p 0mV 3404000p 1mV 3404001p 0mV 3426000p 1mV 3426001p 0mV 3427000p 1mV 3427001p 0mV 3448000p 1mV 3448001p 0mV 3456000p 1mV 3456001p 0mV 3458000p 1mV 3458001p 0mV 3466000p 1mV 3466001p 0mV 3476000p 1mV 3476001p 0mV 3489000p 1mV 3489001p 0mV 3492000p 1mV 3492001p 0mV 3496000p 1mV 3496001p 0mV 3498000p 1mV 3498001p 0mV 3499000p 1mV 3499001p 0mV 3508000p 1mV 3508001p 0mV 3519000p 1mV 3519001p 0mV 3527000p 1mV 3527001p 0mV 3529000p 1mV 3529001p 0mV 3536000p 1mV 3536001p 0mV 3550000p 1mV 3550001p 0mV 3570000p 1mV 3570001p 0mV 3706000p 1mV 3706001p 0mV 3708000p 1mV 3708001p 0mV 3709000p 1mV 3709001p 0mV 3711000p 1mV 3711001p 0mV 3714000p 1mV 3714001p 0mV 3717000p 1mV 3717001p 0mV 3736000p 1mV 3736001p 0mV 3738000p 1mV 3738001p 0mV 3757000p 1mV 3757001p 0mV 3766000p 1mV 3766001p 0mV 3769000p 1mV 3769001p 0mV 3770000p 1mV 3770001p 0mV 3775000p 1mV 3775001p 0mV 3788000p 1mV 3788001p 0mV 3929000p 1mV 3929001p 0mV 3945000p 1mV 3945001p 0mV 3951000p 1mV 3951001p 0mV 3969000p 1mV 3969001p 0mV 3987000p 1mV 3987001p 0mV 3988000p 1mV 3988001p 0mV 3998000p 1mV 3998001p 0mV 4001000p 1mV 4001001p 0mV 4006000p 1mV 4006001p 0mV 4012000p 1mV 4012001p 0mV 4022000p 1mV 4022001p 0mV 4026000p 1mV 4026001p 0mV 4039000p 1mV 4039001p 0mV 4047000p 1mV 4047001p 0mV 4052000p 1mV 4052001p 0mV 4059000p 1mV 4059001p 0mV 4067000p 1mV 4067001p 0mV 4077000p 1mV 4077001p 0mV 4078000p 1mV 4078001p 0mV 4080000p 1mV 4080001p 0mV 4084000p 1mV 4084001p 0mV 4088000p 1mV 4088001p 0mV 4090000p 1mV 4090001p 0mV 4125000p 1mV 4125001p 0mV 4126000p 1mV 4126001p 0mV 4189000p 1mV 4189001p 0mV 4190000p 1mV 4190001p 0mV 4193000p 1mV 4193001p 0mV 4196000p 1mV 4196001p 0mV 4230000p 1mV 4230001p 0mV 4254000p 1mV 4254001p 0mV 4256000p 1mV 4256001p 0mV 4263000p 1mV 4263001p 0mV 4264000p 1mV 4264001p 0mV 4284000p 1mV 4284001p 0mV 4285000p 1mV 4285001p 0mV 4297000p 1mV 4297001p 0mV 4319000p 1mV 4319001p 0mV 4321000p 1mV 4321001p 0mV 4327000p 1mV 4327001p 0mV 4336000p 1mV 4336001p 0mV 4342000p 1mV 4342001p 0mV 4353000p 1mV 4353001p 0mV 4361000p 1mV 4361001p 0mV 4376000p 1mV 4376001p 0mV 4385000p 1mV 4385001p 0mV 4419000p 1mV 4419001p 0mV 4422000p 1mV 4422001p 0mV 4426000p 1mV 4426001p 0mV 4436000p 1mV 4436001p 0mV 4439000p 1mV 4439001p 0mV 4445000p 1mV 4445001p 0mV 4448000p 1mV 4448001p 0mV 4474000p 1mV 4474001p 0mV 4482000p 1mV 4482001p 0mV 4485000p 1mV 4485001p 0mV 4493000p 1mV 4493001p 0mV 4515000p 1mV 4515001p 0mV 4529000p 1mV 4529001p 0mV 4569000p 1mV 4569001p 0mV 4574000p 1mV 4574001p 0mV 4575000p 1mV 4575001p 0mV 4581000p 1mV 4581001p 0mV 4584000p 1mV 4584001p 0mV 4602000p 1mV 4602001p 0mV 4604000p 1mV 4604001p 0mV 4615000p 1mV 4615001p 0mV 4623000p 1mV 4623001p 0mV 4629000p 1mV 4629001p 0mV 4630000p 1mV 4630001p 0mV 4645000p 1mV 4645001p 0mV 4655000p 1mV 4655001p 0mV 4672000p 1mV 4672001p 0mV 4684000p 1mV 4684001p 0mV 4727000p 1mV 4727001p 0mV 4744000p 1mV 4744001p 0mV 4750000p 1mV 4750001p 0mV 4759000p 1mV 4759001p 0mV 4768000p 1mV 4768001p 0mV 4794000p 1mV 4794001p 0mV 4799000p 1mV 4799001p 0mV 4804000p 1mV 4804001p 0mV 4809000p 1mV 4809001p 0mV 4822000p 1mV 4822001p 0mV 4823000p 1mV 4823001p 0mV 4840000p 1mV 4840001p 0mV 4844000p 1mV 4844001p 0mV 4863000p 1mV 4863001p 0mV 4866000p 1mV 4866001p 0mV 4883000p 1mV 4883001p 0mV 4892000p 1mV 4892001p 0mV 4896000p 1mV 4896001p 0mV 4897000p 1mV 4897001p 0mV 4912000p 1mV 4912001p 0mV 4919000p 1mV 4919001p 0mV 4927000p 1mV 4927001p 0mV 4939000p 1mV 4939001p 0mV 4942000p 1mV 4942001p 0mV 4973000p 1mV 4973001p 0mV 4975000p 1mV 4975001p 0mV 4993000p 1mV 4993001p 0mV 5100000p 1mV 5100001p 0mV 5107000p 1mV 5107001p 0mV 5125000p 1mV 5125001p 0mV 5130000p 1mV 5130001p 0mV 5134000p 1mV 5134001p 0mV 5140000p 1mV 5140001p 0mV 5142000p 1mV 5142001p 0mV 5146000p 1mV 5146001p 0mV 5164000p 1mV 5164001p 0mV 5166000p 1mV 5166001p 0mV 5175000p 1mV 5175001p 0mV 5203000p 1mV 5203001p 0mV 5207000p 1mV 5207001p 0mV 5217000p 1mV 5217001p 0mV 5232000p 1mV 5232001p 0mV 5233000p 1mV 5233001p 0mV 5238000p 1mV 5238001p 0mV 5241000p 1mV 5241001p 0mV 5255000p 1mV 5255001p 0mV 5267000p 1mV 5267001p 0mV 5269000p 1mV 5269001p 0mV 5282000p 1mV 5282001p 0mV 5284000p 1mV 5284001p 0mV 5298000p 1mV 5298001p 0mV 5310000p 1mV 5310001p 0mV 5326000p 1mV 5326001p 0mV 5328000p 1mV 5328001p 0mV 5351000p 1mV 5351001p 0mV 5361000p 1mV 5361001p 0mV 5364000p 1mV 5364001p 0mV 5389000p 1mV 5389001p 0mV 5916000p 1mV 5916001p 0mV 5931000p 1mV 5931001p 0mV 5936000p 1mV 5936001p 0mV 5939000p 1mV 5939001p 0mV 5955000p 1mV 5955001p 0mV 5965000p 1mV 5965001p 0mV 5966000p 1mV 5966001p 0mV 5972000p 1mV 5972001p 0mV 5979000p 1mV 5979001p 0mV 6100000p 1mV 6100001p 0mV 6115000p 1mV 6115001p 0mV 6116000p 1mV 6116001p 0mV 6126000p 1mV 6126001p 0mV 6172000p 1mV 6172001p 0mV 6183000p 1mV 6183001p 0mV 6192000p 1mV 6192001p 0mV 6701000p 1mV 6701001p 0mV 6723000p 1mV 6723001p 0mV 6725000p 1mV 6725001p 0mV 6741000p 1mV 6741001p 0mV 6745000p 1mV 6745001p 0mV 6754000p 1mV 6754001p 0mV 6762000p 1mV 6762001p 0mV 6792000p 1mV 6792001p 0mV 6814000p 1mV 6814001p 0mV 6822000p 1mV 6822001p 0mV 6825000p 1mV 6825001p 0mV 6835000p 1mV 6835001p 0mV 6838000p 1mV 6838001p 0mV 6859000p 1mV 6859001p 0mV 6866000p 1mV 6866001p 0mV 6870000p 1mV 6870001p 0mV 6877000p 1mV 6877001p 0mV 6888000p 1mV 6888001p 0mV 6894000p 1mV 6894001p 0mV 7174000p 1mV 7174001p 0mV 7309000p 1mV 7309001p 0mV 7372000p 1mV 7372001p 0mV 7376000p 1mV 7376001p 0mV 7742000p 1mV 7742001p 0mV 8825000p 1mV 8825001p 0mV 8829000p 1mV 8829001p 0mV 8840000p 1mV 8840001p 0mV 8847000p 1mV 8847001p 0mV 8849000p 1mV 8849001p 0mV 8884000p 1mV 8884001p 0mV 8886000p 1mV 8886001p 0mV 9619000p 1mV 9619001p 0mV 9634000p 1mV 9634001p 0mV 9648000p 1mV 9648001p 0mV 9687000p 1mV 9687001p 0mV 9696000p 1mV 9696001p 0mV 9699000p 1mV 9699001p 0mV 9712000p 1mV 9712001p 0mV 9734000p 1mV 9734001p 0mV 9745000p 1mV 9745001p 0mV 9757000p 1mV 9757001p 0mV 9758000p 1mV 9758001p 0mV 9761000p 1mV 9761001p 0mV 9780000p 1mV 9780001p 0mV 9798000p 1mV 9798001p 0mV 9806000p 1mV 9806001p 0mV 9808000p 1mV 9808001p 0mV 9824000p 1mV 9824001p 0mV 9830000p 1mV 9830001p 0mV 9831000p 1mV 9831001p 0mV 9838000p 1mV 9838001p 0mV 9846000p 1mV 9846001p 0mV 9857000p 1mV 9857001p 0mV 9861000p 1mV 9861001p 0mV 9865000p 1mV 9865001p 0mV 9870000p 1mV 9870001p 0mV 9872000p 1mV 9872001p 0mV 9877000p 1mV 9877001p 0mV 9882000p 1mV 9882001p 0mV 9892000p 1mV 9892001p 0mV 9915000p 1mV 9915001p 0mV 9916000p 1mV 9916001p 0mV 9919000p 1mV 9919001p 0mV 9944000p 1mV 9944001p 0mV 9956000p 1mV 9956001p 0mV 9957000p 1mV 9957001p 0mV 9962000p 1mV 9962001p 0mV 9973000p 1mV 9973001p 0mV 9984000p 1mV 9984001p 0mV 9991000p 1mV 9991001p 0mV 9993000p 1mV 9993001p 0mV 9994000p 1mV 9994001p 0mV)
.ENDS conductors__anyBias-Lk_0_702

.SUBCKT conductors__anyBias-Lk_0_703 bottom out
VrampSppl@0 bottom out pwl (100000p 1mV 100001p 0mV 101000p 1mV 101001p 0mV 130000p 1mV 130001p 0mV 177000p 1mV 177001p 0mV 302000p 1mV 302001p 0mV 303000p 1mV 303001p 0mV 316000p 1mV 316001p 0mV 333000p 1mV 333001p 0mV 339000p 1mV 339001p 0mV 343000p 1mV 343001p 0mV 346000p 1mV 346001p 0mV 349000p 1mV 349001p 0mV 352000p 1mV 352001p 0mV 358000p 1mV 358001p 0mV 375000p 1mV 375001p 0mV 391000p 1mV 391001p 0mV 394000p 1mV 394001p 0mV 405000p 1mV 405001p 0mV 430000p 1mV 430001p 0mV 432000p 1mV 432001p 0mV 475000p 1mV 475001p 0mV 499000p 1mV 499001p 0mV 504000p 1mV 504001p 0mV 525000p 1mV 525001p 0mV 527000p 1mV 527001p 0mV 535000p 1mV 535001p 0mV 539000p 1mV 539001p 0mV 563000p 1mV 563001p 0mV 614000p 1mV 614001p 0mV 633000p 1mV 633001p 0mV 641000p 1mV 641001p 0mV 716000p 1mV 716001p 0mV 718000p 1mV 718001p 0mV 729000p 1mV 729001p 0mV 739000p 1mV 739001p 0mV 741000p 1mV 741001p 0mV 749000p 1mV 749001p 0mV 757000p 1mV 757001p 0mV 767000p 1mV 767001p 0mV 810000p 1mV 810001p 0mV 850000p 1mV 850001p 0mV 856000p 1mV 856001p 0mV 867000p 1mV 867001p 0mV 898000p 1mV 898001p 0mV 906000p 1mV 906001p 0mV 919000p 1mV 919001p 0mV 941000p 1mV 941001p 0mV 945000p 1mV 945001p 0mV 946000p 1mV 946001p 0mV 971000p 1mV 971001p 0mV 973000p 1mV 973001p 0mV 1034000p 1mV 1034001p 0mV 1044000p 1mV 1044001p 0mV 1050000p 1mV 1050001p 0mV 1067000p 1mV 1067001p 0mV 1083000p 1mV 1083001p 0mV 1095000p 1mV 1095001p 0mV 1096000p 1mV 1096001p 0mV 1112000p 1mV 1112001p 0mV 1114000p 1mV 1114001p 0mV 1117000p 1mV 1117001p 0mV 1119000p 1mV 1119001p 0mV 1136000p 1mV 1136001p 0mV 1151000p 1mV 1151001p 0mV 1152000p 1mV 1152001p 0mV 1162000p 1mV 1162001p 0mV 1169000p 1mV 1169001p 0mV 1182000p 1mV 1182001p 0mV 1201000p 1mV 1201001p 0mV 1221000p 1mV 1221001p 0mV 1248000p 1mV 1248001p 0mV 1258000p 1mV 1258001p 0mV 1280000p 1mV 1280001p 0mV 1282000p 1mV 1282001p 0mV 1302000p 1mV 1302001p 0mV 1304000p 1mV 1304001p 0mV 1333000p 1mV 1333001p 0mV 1336000p 1mV 1336001p 0mV 1344000p 1mV 1344001p 0mV 1397000p 1mV 1397001p 0mV 1436000p 1mV 1436001p 0mV 1449000p 1mV 1449001p 0mV 1470000p 1mV 1470001p 0mV 1477000p 1mV 1477001p 0mV 1489000p 1mV 1489001p 0mV 1523000p 1mV 1523001p 0mV 1524000p 1mV 1524001p 0mV 1526000p 1mV 1526001p 0mV 1553000p 1mV 1553001p 0mV 1563000p 1mV 1563001p 0mV 1568000p 1mV 1568001p 0mV 1570000p 1mV 1570001p 0mV 1571000p 1mV 1571001p 0mV 1589000p 1mV 1589001p 0mV 1603000p 1mV 1603001p 0mV 1618000p 1mV 1618001p 0mV 1621000p 1mV 1621001p 0mV 1626000p 1mV 1626001p 0mV 1688000p 1mV 1688001p 0mV 1691000p 1mV 1691001p 0mV 1700000p 1mV 1700001p 0mV 1724000p 1mV 1724001p 0mV 1772000p 1mV 1772001p 0mV 1779000p 1mV 1779001p 0mV 1790000p 1mV 1790001p 0mV 1798000p 1mV 1798001p 0mV 1807000p 1mV 1807001p 0mV 1808000p 1mV 1808001p 0mV 1811000p 1mV 1811001p 0mV 1815000p 1mV 1815001p 0mV 1820000p 1mV 1820001p 0mV 1833000p 1mV 1833001p 0mV 1837000p 1mV 1837001p 0mV 1861000p 1mV 1861001p 0mV 1873000p 1mV 1873001p 0mV 1882000p 1mV 1882001p 0mV 1910000p 1mV 1910001p 0mV 1919000p 1mV 1919001p 0mV 1959000p 1mV 1959001p 0mV 1986000p 1mV 1986001p 0mV 1994000p 1mV 1994001p 0mV 2038000p 1mV 2038001p 0mV 2049000p 1mV 2049001p 0mV 2053000p 1mV 2053001p 0mV 2054000p 1mV 2054001p 0mV 2055000p 1mV 2055001p 0mV 2058000p 1mV 2058001p 0mV 2068000p 1mV 2068001p 0mV 2080000p 1mV 2080001p 0mV 2089000p 1mV 2089001p 0mV 2096000p 1mV 2096001p 0mV 2108000p 1mV 2108001p 0mV 2119000p 1mV 2119001p 0mV 2137000p 1mV 2137001p 0mV 2140000p 1mV 2140001p 0mV 2157000p 1mV 2157001p 0mV 2158000p 1mV 2158001p 0mV 2180000p 1mV 2180001p 0mV 2196000p 1mV 2196001p 0mV 2207000p 1mV 2207001p 0mV 2226000p 1mV 2226001p 0mV 2245000p 1mV 2245001p 0mV 2290000p 1mV 2290001p 0mV 2309000p 1mV 2309001p 0mV 2376000p 1mV 2376001p 0mV 2382000p 1mV 2382001p 0mV 2384000p 1mV 2384001p 0mV 2402000p 1mV 2402001p 0mV 2405000p 1mV 2405001p 0mV 2411000p 1mV 2411001p 0mV 2436000p 1mV 2436001p 0mV 2440000p 1mV 2440001p 0mV 2449000p 1mV 2449001p 0mV 2452000p 1mV 2452001p 0mV 2524000p 1mV 2524001p 0mV 2532000p 1mV 2532001p 0mV 2539000p 1mV 2539001p 0mV 2544000p 1mV 2544001p 0mV 2548000p 1mV 2548001p 0mV 2551000p 1mV 2551001p 0mV 2552000p 1mV 2552001p 0mV 2589000p 1mV 2589001p 0mV 2593000p 1mV 2593001p 0mV 2594000p 1mV 2594001p 0mV 2601000p 1mV 2601001p 0mV 2603000p 1mV 2603001p 0mV 2629000p 1mV 2629001p 0mV 2630000p 1mV 2630001p 0mV 2636000p 1mV 2636001p 0mV 2643000p 1mV 2643001p 0mV 2658000p 1mV 2658001p 0mV 2665000p 1mV 2665001p 0mV 2672000p 1mV 2672001p 0mV 2682000p 1mV 2682001p 0mV 2686000p 1mV 2686001p 0mV 2693000p 1mV 2693001p 0mV 2695000p 1mV 2695001p 0mV 2697000p 1mV 2697001p 0mV 2698000p 1mV 2698001p 0mV 2708000p 1mV 2708001p 0mV 2747000p 1mV 2747001p 0mV 2755000p 1mV 2755001p 0mV 2787000p 1mV 2787001p 0mV 2794000p 1mV 2794001p 0mV 2796000p 1mV 2796001p 0mV 2803000p 1mV 2803001p 0mV 2811000p 1mV 2811001p 0mV 2824000p 1mV 2824001p 0mV 2848000p 1mV 2848001p 0mV 2865000p 1mV 2865001p 0mV 2870000p 1mV 2870001p 0mV 2872000p 1mV 2872001p 0mV 2883000p 1mV 2883001p 0mV 2889000p 1mV 2889001p 0mV 2894000p 1mV 2894001p 0mV 2918000p 1mV 2918001p 0mV 2926000p 1mV 2926001p 0mV 2939000p 1mV 2939001p 0mV 2969000p 1mV 2969001p 0mV 3000000p 1mV 3000001p 0mV 3039000p 1mV 3039001p 0mV 3070000p 1mV 3070001p 0mV 3077000p 1mV 3077001p 0mV 3078000p 1mV 3078001p 0mV 3111000p 1mV 3111001p 0mV 3122000p 1mV 3122001p 0mV 3126000p 1mV 3126001p 0mV 3127000p 1mV 3127001p 0mV 3129000p 1mV 3129001p 0mV 3141000p 1mV 3141001p 0mV 3155000p 1mV 3155001p 0mV 3167000p 1mV 3167001p 0mV 3189000p 1mV 3189001p 0mV 3206000p 1mV 3206001p 0mV 3219000p 1mV 3219001p 0mV 3234000p 1mV 3234001p 0mV 3249000p 1mV 3249001p 0mV 3254000p 1mV 3254001p 0mV 3263000p 1mV 3263001p 0mV 3264000p 1mV 3264001p 0mV 3270000p 1mV 3270001p 0mV 3300000p 1mV 3300001p 0mV 3301000p 1mV 3301001p 0mV 3303000p 1mV 3303001p 0mV 3384000p 1mV 3384001p 0mV 3395000p 1mV 3395001p 0mV 3409000p 1mV 3409001p 0mV 3418000p 1mV 3418001p 0mV 3425000p 1mV 3425001p 0mV 3454000p 1mV 3454001p 0mV 3462000p 1mV 3462001p 0mV 3469000p 1mV 3469001p 0mV 3476000p 1mV 3476001p 0mV 3495000p 1mV 3495001p 0mV 3498000p 1mV 3498001p 0mV 3502000p 1mV 3502001p 0mV 3503000p 1mV 3503001p 0mV 3527000p 1mV 3527001p 0mV 3537000p 1mV 3537001p 0mV 3544000p 1mV 3544001p 0mV 3553000p 1mV 3553001p 0mV 3565000p 1mV 3565001p 0mV 3574000p 1mV 3574001p 0mV 3598000p 1mV 3598001p 0mV 3663000p 1mV 3663001p 0mV 3700000p 1mV 3700001p 0mV 3701000p 1mV 3701001p 0mV 3755000p 1mV 3755001p 0mV 3770000p 1mV 3770001p 0mV 3779000p 1mV 3779001p 0mV 3780000p 1mV 3780001p 0mV 3836000p 1mV 3836001p 0mV 3842000p 1mV 3842001p 0mV 3856000p 1mV 3856001p 0mV 3920000p 1mV 3920001p 0mV 3921000p 1mV 3921001p 0mV 3933000p 1mV 3933001p 0mV 3947000p 1mV 3947001p 0mV 3957000p 1mV 3957001p 0mV 3964000p 1mV 3964001p 0mV 4000000p 1mV 4000001p 0mV 4006000p 1mV 4006001p 0mV 4043000p 1mV 4043001p 0mV 4051000p 1mV 4051001p 0mV 4057000p 1mV 4057001p 0mV 4075000p 1mV 4075001p 0mV 4080000p 1mV 4080001p 0mV 4097000p 1mV 4097001p 0mV 4102000p 1mV 4102001p 0mV 4118000p 1mV 4118001p 0mV 4129000p 1mV 4129001p 0mV 4146000p 1mV 4146001p 0mV 4187000p 1mV 4187001p 0mV 4218000p 1mV 4218001p 0mV 4232000p 1mV 4232001p 0mV 4241000p 1mV 4241001p 0mV 4316000p 1mV 4316001p 0mV 4319000p 1mV 4319001p 0mV 4349000p 1mV 4349001p 0mV 4421000p 1mV 4421001p 0mV 4446000p 1mV 4446001p 0mV 4454000p 1mV 4454001p 0mV 4465000p 1mV 4465001p 0mV 4471000p 1mV 4471001p 0mV 4478000p 1mV 4478001p 0mV 4554000p 1mV 4554001p 0mV 4577000p 1mV 4577001p 0mV 4606000p 1mV 4606001p 0mV 4611000p 1mV 4611001p 0mV 4643000p 1mV 4643001p 0mV 4661000p 1mV 4661001p 0mV 4672000p 1mV 4672001p 0mV 4688000p 1mV 4688001p 0mV 4693000p 1mV 4693001p 0mV 4720000p 1mV 4720001p 0mV 4731000p 1mV 4731001p 0mV 4734000p 1mV 4734001p 0mV 4737000p 1mV 4737001p 0mV 4804000p 1mV 4804001p 0mV 4806000p 1mV 4806001p 0mV 4877000p 1mV 4877001p 0mV 4891000p 1mV 4891001p 0mV 4975000p 1mV 4975001p 0mV 4977000p 1mV 4977001p 0mV 5033000p 1mV 5033001p 0mV 5070000p 1mV 5070001p 0mV 5090000p 1mV 5090001p 0mV 5095000p 1mV 5095001p 0mV 5114000p 1mV 5114001p 0mV 5119000p 1mV 5119001p 0mV 5128000p 1mV 5128001p 0mV 5136000p 1mV 5136001p 0mV 5138000p 1mV 5138001p 0mV 5155000p 1mV 5155001p 0mV 5176000p 1mV 5176001p 0mV 5178000p 1mV 5178001p 0mV 5201000p 1mV 5201001p 0mV 5211000p 1mV 5211001p 0mV 5221000p 1mV 5221001p 0mV 5244000p 1mV 5244001p 0mV 5275000p 1mV 5275001p 0mV 5308000p 1mV 5308001p 0mV 5309000p 1mV 5309001p 0mV 5328000p 1mV 5328001p 0mV 5393000p 1mV 5393001p 0mV 5485000p 1mV 5485001p 0mV 5575000p 1mV 5575001p 0mV 5601000p 1mV 5601001p 0mV 5649000p 1mV 5649001p 0mV 5660000p 1mV 5660001p 0mV 5661000p 1mV 5661001p 0mV 5665000p 1mV 5665001p 0mV 5683000p 1mV 5683001p 0mV 5758000p 1mV 5758001p 0mV 5774000p 1mV 5774001p 0mV 5806000p 1mV 5806001p 0mV 5835000p 1mV 5835001p 0mV 5857000p 1mV 5857001p 0mV 5940000p 1mV 5940001p 0mV 5944000p 1mV 5944001p 0mV 5963000p 1mV 5963001p 0mV 5965000p 1mV 5965001p 0mV 5967000p 1mV 5967001p 0mV 5974000p 1mV 5974001p 0mV 5987000p 1mV 5987001p 0mV 5992000p 1mV 5992001p 0mV 6031000p 1mV 6031001p 0mV 6083000p 1mV 6083001p 0mV 6094000p 1mV 6094001p 0mV 6103000p 1mV 6103001p 0mV 6106000p 1mV 6106001p 0mV 6115000p 1mV 6115001p 0mV 6116000p 1mV 6116001p 0mV 6119000p 1mV 6119001p 0mV 6139000p 1mV 6139001p 0mV 6153000p 1mV 6153001p 0mV 6163000p 1mV 6163001p 0mV 6170000p 1mV 6170001p 0mV 6181000p 1mV 6181001p 0mV 6220000p 1mV 6220001p 0mV 6246000p 1mV 6246001p 0mV 6250000p 1mV 6250001p 0mV 6261000p 1mV 6261001p 0mV 6267000p 1mV 6267001p 0mV 6275000p 1mV 6275001p 0mV 6295000p 1mV 6295001p 0mV 6298000p 1mV 6298001p 0mV 6321000p 1mV 6321001p 0mV 6330000p 1mV 6330001p 0mV 6356000p 1mV 6356001p 0mV 6370000p 1mV 6370001p 0mV 6372000p 1mV 6372001p 0mV 6438000p 1mV 6438001p 0mV 6439000p 1mV 6439001p 0mV 6442000p 1mV 6442001p 0mV 6456000p 1mV 6456001p 0mV 6458000p 1mV 6458001p 0mV 6481000p 1mV 6481001p 0mV 6499000p 1mV 6499001p 0mV 6517000p 1mV 6517001p 0mV 6538000p 1mV 6538001p 0mV 6554000p 1mV 6554001p 0mV 6562000p 1mV 6562001p 0mV 6563000p 1mV 6563001p 0mV 6624000p 1mV 6624001p 0mV 6685000p 1mV 6685001p 0mV 6698000p 1mV 6698001p 0mV 6705000p 1mV 6705001p 0mV 6706000p 1mV 6706001p 0mV 6711000p 1mV 6711001p 0mV 6715000p 1mV 6715001p 0mV 6721000p 1mV 6721001p 0mV 6758000p 1mV 6758001p 0mV 6759000p 1mV 6759001p 0mV 6766000p 1mV 6766001p 0mV 6783000p 1mV 6783001p 0mV 6785000p 1mV 6785001p 0mV 6849000p 1mV 6849001p 0mV 6869000p 1mV 6869001p 0mV 6883000p 1mV 6883001p 0mV 6905000p 1mV 6905001p 0mV 6906000p 1mV 6906001p 0mV 6933000p 1mV 6933001p 0mV 6948000p 1mV 6948001p 0mV 6958000p 1mV 6958001p 0mV 6962000p 1mV 6962001p 0mV 6998000p 1mV 6998001p 0mV 7011000p 1mV 7011001p 0mV 7078000p 1mV 7078001p 0mV 7084000p 1mV 7084001p 0mV 7093000p 1mV 7093001p 0mV 7105000p 1mV 7105001p 0mV 7120000p 1mV 7120001p 0mV 7175000p 1mV 7175001p 0mV 7182000p 1mV 7182001p 0mV 7262000p 1mV 7262001p 0mV 7263000p 1mV 7263001p 0mV 7284000p 1mV 7284001p 0mV 7289000p 1mV 7289001p 0mV 7311000p 1mV 7311001p 0mV 7317000p 1mV 7317001p 0mV 7323000p 1mV 7323001p 0mV 7331000p 1mV 7331001p 0mV 7332000p 1mV 7332001p 0mV 7355000p 1mV 7355001p 0mV 7359000p 1mV 7359001p 0mV 7362000p 1mV 7362001p 0mV 7392000p 1mV 7392001p 0mV 7397000p 1mV 7397001p 0mV 7488000p 1mV 7488001p 0mV 7524000p 1mV 7524001p 0mV 7534000p 1mV 7534001p 0mV 7548000p 1mV 7548001p 0mV 7573000p 1mV 7573001p 0mV 7579000p 1mV 7579001p 0mV 7617000p 1mV 7617001p 0mV 7632000p 1mV 7632001p 0mV 7698000p 1mV 7698001p 0mV 7730000p 1mV 7730001p 0mV 7746000p 1mV 7746001p 0mV 7754000p 1mV 7754001p 0mV 7763000p 1mV 7763001p 0mV 7770000p 1mV 7770001p 0mV 7778000p 1mV 7778001p 0mV 7782000p 1mV 7782001p 0mV 7785000p 1mV 7785001p 0mV 7855000p 1mV 7855001p 0mV 7872000p 1mV 7872001p 0mV 7876000p 1mV 7876001p 0mV 7889000p 1mV 7889001p 0mV 7909000p 1mV 7909001p 0mV 7911000p 1mV 7911001p 0mV 7960000p 1mV 7960001p 0mV 7965000p 1mV 7965001p 0mV 7966000p 1mV 7966001p 0mV 7990000p 1mV 7990001p 0mV 8000000p 1mV 8000001p 0mV 8012000p 1mV 8012001p 0mV 8049000p 1mV 8049001p 0mV 8062000p 1mV 8062001p 0mV 8064000p 1mV 8064001p 0mV 8072000p 1mV 8072001p 0mV 8087000p 1mV 8087001p 0mV 8106000p 1mV 8106001p 0mV 8111000p 1mV 8111001p 0mV 8136000p 1mV 8136001p 0mV 8149000p 1mV 8149001p 0mV 8209000p 1mV 8209001p 0mV 8259000p 1mV 8259001p 0mV 8262000p 1mV 8262001p 0mV 8267000p 1mV 8267001p 0mV 8296000p 1mV 8296001p 0mV 8300000p 1mV 8300001p 0mV 8301000p 1mV 8301001p 0mV 8306000p 1mV 8306001p 0mV 8314000p 1mV 8314001p 0mV 8345000p 1mV 8345001p 0mV 8378000p 1mV 8378001p 0mV 8380000p 1mV 8380001p 0mV 8385000p 1mV 8385001p 0mV 8434000p 1mV 8434001p 0mV 8442000p 1mV 8442001p 0mV 8449000p 1mV 8449001p 0mV 8482000p 1mV 8482001p 0mV 8501000p 1mV 8501001p 0mV 8505000p 1mV 8505001p 0mV 8521000p 1mV 8521001p 0mV 8526000p 1mV 8526001p 0mV 8532000p 1mV 8532001p 0mV 8559000p 1mV 8559001p 0mV 8574000p 1mV 8574001p 0mV 8580000p 1mV 8580001p 0mV 8608000p 1mV 8608001p 0mV 8609000p 1mV 8609001p 0mV 8638000p 1mV 8638001p 0mV 8645000p 1mV 8645001p 0mV 8653000p 1mV 8653001p 0mV 8669000p 1mV 8669001p 0mV 8670000p 1mV 8670001p 0mV 8674000p 1mV 8674001p 0mV 8683000p 1mV 8683001p 0mV 8728000p 1mV 8728001p 0mV 8759000p 1mV 8759001p 0mV 8767000p 1mV 8767001p 0mV 8772000p 1mV 8772001p 0mV 8790000p 1mV 8790001p 0mV 8802000p 1mV 8802001p 0mV 8807000p 1mV 8807001p 0mV 8812000p 1mV 8812001p 0mV 8815000p 1mV 8815001p 0mV 8818000p 1mV 8818001p 0mV 8825000p 1mV 8825001p 0mV 8863000p 1mV 8863001p 0mV 8883000p 1mV 8883001p 0mV 8884000p 1mV 8884001p 0mV 8891000p 1mV 8891001p 0mV 8897000p 1mV 8897001p 0mV 8944000p 1mV 8944001p 0mV 8946000p 1mV 8946001p 0mV 8976000p 1mV 8976001p 0mV 8992000p 1mV 8992001p 0mV 8995000p 1mV 8995001p 0mV 9008000p 1mV 9008001p 0mV 9021000p 1mV 9021001p 0mV 9061000p 1mV 9061001p 0mV 9114000p 1mV 9114001p 0mV 9185000p 1mV 9185001p 0mV 9197000p 1mV 9197001p 0mV 9239000p 1mV 9239001p 0mV 9280000p 1mV 9280001p 0mV 9288000p 1mV 9288001p 0mV 9302000p 1mV 9302001p 0mV 9324000p 1mV 9324001p 0mV 9333000p 1mV 9333001p 0mV 9335000p 1mV 9335001p 0mV 9342000p 1mV 9342001p 0mV 9369000p 1mV 9369001p 0mV 9373000p 1mV 9373001p 0mV 9375000p 1mV 9375001p 0mV 9380000p 1mV 9380001p 0mV 9394000p 1mV 9394001p 0mV 9422000p 1mV 9422001p 0mV 9425000p 1mV 9425001p 0mV 9426000p 1mV 9426001p 0mV 9428000p 1mV 9428001p 0mV 9445000p 1mV 9445001p 0mV 9459000p 1mV 9459001p 0mV 9465000p 1mV 9465001p 0mV 9474000p 1mV 9474001p 0mV 9493000p 1mV 9493001p 0mV 9505000p 1mV 9505001p 0mV 9550000p 1mV 9550001p 0mV 9575000p 1mV 9575001p 0mV 9581000p 1mV 9581001p 0mV 9589000p 1mV 9589001p 0mV 9594000p 1mV 9594001p 0mV 9610000p 1mV 9610001p 0mV 9631000p 1mV 9631001p 0mV 9644000p 1mV 9644001p 0mV 9686000p 1mV 9686001p 0mV 9713000p 1mV 9713001p 0mV 9767000p 1mV 9767001p 0mV 9769000p 1mV 9769001p 0mV 9770000p 1mV 9770001p 0mV 9799000p 1mV 9799001p 0mV 9802000p 1mV 9802001p 0mV 9816000p 1mV 9816001p 0mV 9853000p 1mV 9853001p 0mV 9854000p 1mV 9854001p 0mV 9861000p 1mV 9861001p 0mV 9876000p 1mV 9876001p 0mV 9886000p 1mV 9886001p 0mV 9889000p 1mV 9889001p 0mV 9893000p 1mV 9893001p 0mV 9919000p 1mV 9919001p 0mV 9998000p 1mV 9998001p 0mV)
.ENDS conductors__anyBias-Lk_0_703

.SUBCKT conductors__anyBias-Lk_0_704 bottom out
VrampSppl@0 bottom out pwl(0p 1mV 1p 0mV 12000p 1mV 12001p 0mV 15000p 1mV 15001p 0mV 17000p 1mV 17001p 0mV 20000p 1mV 20001p 0mV 34000p 1mV 34001p 0mV 35000p 1mV 35001p 0mV 40000p 1mV 40001p 0mV 46000p 1mV 46001p 0mV 58000p 1mV 58001p 0mV 67000p 1mV 67001p 0mV 70000p 1mV 70001p 0mV 93000p 1mV 93001p 0mV 125000p 1mV 125001p 0mV 127000p 1mV 127001p 0mV 129000p 1mV 129001p 0mV 138000p 1mV 138001p 0mV 170000p 1mV 170001p 0mV 175000p 1mV 175001p 0mV 180000p 1mV 180001p 0mV 190000p 1mV 190001p 0mV 196000p 1mV 196001p 0mV 200000p 1mV 200001p 0mV 210000p 1mV 210001p 0mV 211000p 1mV 211001p 0mV 251000p 1mV 251001p 0mV 284000p 1mV 284001p 0mV 287000p 1mV 287001p 0mV 288000p 1mV 288001p 0mV 290000p 1mV 290001p 0mV 297000p 1mV 297001p 0mV 299000p 1mV 299001p 0mV 1604000p 1mV 1604001p 0mV 1606000p 1mV 1606001p 0mV 1609000p 1mV 1609001p 0mV 1613000p 1mV 1613001p 0mV 1624000p 1mV 1624001p 0mV 1628000p 1mV 1628001p 0mV 1652000p 1mV 1652001p 0mV 1654000p 1mV 1654001p 0mV 1657000p 1mV 1657001p 0mV 1672000p 1mV 1672001p 0mV 1687000p 1mV 1687001p 0mV 1689000p 1mV 1689001p 0mV 1814000p 1mV 1814001p 0mV 1819000p 1mV 1819001p 0mV 1824000p 1mV 1824001p 0mV 1825000p 1mV 1825001p 0mV 1827000p 1mV 1827001p 0mV 1840000p 1mV 1840001p 0mV 1864000p 1mV 1864001p 0mV 1875000p 1mV 1875001p 0mV 1883000p 1mV 1883001p 0mV 2001000p 1mV 2001001p 0mV 2023000p 1mV 2023001p 0mV 2035000p 1mV 2035001p 0mV 2042000p 1mV 2042001p 0mV 2049000p 1mV 2049001p 0mV 2057000p 1mV 2057001p 0mV 2068000p 1mV 2068001p 0mV 2076000p 1mV 2076001p 0mV 2078000p 1mV 2078001p 0mV 2087000p 1mV 2087001p 0mV 2208000p 1mV 2208001p 0mV 2211000p 1mV 2211001p 0mV 2213000p 1mV 2213001p 0mV 2221000p 1mV 2221001p 0mV 2228000p 1mV 2228001p 0mV 2236000p 1mV 2236001p 0mV 2248000p 1mV 2248001p 0mV 2258000p 1mV 2258001p 0mV 2264000p 1mV 2264001p 0mV 2275000p 1mV 2275001p 0mV 2288000p 1mV 2288001p 0mV 2301000p 1mV 2301001p 0mV 2302000p 1mV 2302001p 0mV 2316000p 1mV 2316001p 0mV 2332000p 1mV 2332001p 0mV 2357000p 1mV 2357001p 0mV 2360000p 1mV 2360001p 0mV 2368000p 1mV 2368001p 0mV 2374000p 1mV 2374001p 0mV 2390000p 1mV 2390001p 0mV 2401000p 1mV 2401001p 0mV 2408000p 1mV 2408001p 0mV 2417000p 1mV 2417001p 0mV 2441000p 1mV 2441001p 0mV 2451000p 1mV 2451001p 0mV 2456000p 1mV 2456001p 0mV 2489000p 1mV 2489001p 0mV 2492000p 1mV 2492001p 0mV 2494000p 1mV 2494001p 0mV 2495000p 1mV 2495001p 0mV 2506000p 1mV 2506001p 0mV 2509000p 1mV 2509001p 0mV 2523000p 1mV 2523001p 0mV 2524000p 1mV 2524001p 0mV 2529000p 1mV 2529001p 0mV 2530000p 1mV 2530001p 0mV 2547000p 1mV 2547001p 0mV 2550000p 1mV 2550001p 0mV 2556000p 1mV 2556001p 0mV 2559000p 1mV 2559001p 0mV 2561000p 1mV 2561001p 0mV 2565000p 1mV 2565001p 0mV 2577000p 1mV 2577001p 0mV 2582000p 1mV 2582001p 0mV 2587000p 1mV 2587001p 0mV 2594000p 1mV 2594001p 0mV 2600000p 1mV 2600001p 0mV 2610000p 1mV 2610001p 0mV 2622000p 1mV 2622001p 0mV 2626000p 1mV 2626001p 0mV 2641000p 1mV 2641001p 0mV 2646000p 1mV 2646001p 0mV 2657000p 1mV 2657001p 0mV 2663000p 1mV 2663001p 0mV 2678000p 1mV 2678001p 0mV 2691000p 1mV 2691001p 0mV 2693000p 1mV 2693001p 0mV 2697000p 1mV 2697001p 0mV 2707000p 1mV 2707001p 0mV 2712000p 1mV 2712001p 0mV 2713000p 1mV 2713001p 0mV 2721000p 1mV 2721001p 0mV 2729000p 1mV 2729001p 0mV 2743000p 1mV 2743001p 0mV 2758000p 1mV 2758001p 0mV 2770000p 1mV 2770001p 0mV 2772000p 1mV 2772001p 0mV 2779000p 1mV 2779001p 0mV 2811000p 1mV 2811001p 0mV 2812000p 1mV 2812001p 0mV 2817000p 1mV 2817001p 0mV 2821000p 1mV 2821001p 0mV 2823000p 1mV 2823001p 0mV 2827000p 1mV 2827001p 0mV 2832000p 1mV 2832001p 0mV 2844000p 1mV 2844001p 0mV 2852000p 1mV 2852001p 0mV 2861000p 1mV 2861001p 0mV 2863000p 1mV 2863001p 0mV 2866000p 1mV 2866001p 0mV 2875000p 1mV 2875001p 0mV 2877000p 1mV 2877001p 0mV 2878000p 1mV 2878001p 0mV 2882000p 1mV 2882001p 0mV 2884000p 1mV 2884001p 0mV 2892000p 1mV 2892001p 0mV 2902000p 1mV 2902001p 0mV 2922000p 1mV 2922001p 0mV 2929000p 1mV 2929001p 0mV 2931000p 1mV 2931001p 0mV 2934000p 1mV 2934001p 0mV 2969000p 1mV 2969001p 0mV 2971000p 1mV 2971001p 0mV 2982000p 1mV 2982001p 0mV 2983000p 1mV 2983001p 0mV 2993000p 1mV 2993001p 0mV 3005000p 1mV 3005001p 0mV 3006000p 1mV 3006001p 0mV 3010000p 1mV 3010001p 0mV 3029000p 1mV 3029001p 0mV 3031000p 1mV 3031001p 0mV 3034000p 1mV 3034001p 0mV 3047000p 1mV 3047001p 0mV 3052000p 1mV 3052001p 0mV 3063000p 1mV 3063001p 0mV 3085000p 1mV 3085001p 0mV 3090000p 1mV 3090001p 0mV 3600000p 1mV 3600001p 0mV 3608000p 1mV 3608001p 0mV 3609000p 1mV 3609001p 0mV 3610000p 1mV 3610001p 0mV 3629000p 1mV 3629001p 0mV 3643000p 1mV 3643001p 0mV 3659000p 1mV 3659001p 0mV 3660000p 1mV 3660001p 0mV 3815000p 1mV 3815001p 0mV 3821000p 1mV 3821001p 0mV 3839000p 1mV 3839001p 0mV 3856000p 1mV 3856001p 0mV 3868000p 1mV 3868001p 0mV 3884000p 1mV 3884001p 0mV 3897000p 1mV 3897001p 0mV 5007000p 1mV 5007001p 0mV 5008000p 1mV 5008001p 0mV 5013000p 1mV 5013001p 0mV 5015000p 1mV 5015001p 0mV 5019000p 1mV 5019001p 0mV 5020000p 1mV 5020001p 0mV 5053000p 1mV 5053001p 0mV 5064000p 1mV 5064001p 0mV 5066000p 1mV 5066001p 0mV 5082000p 1mV 5082001p 0mV 5093000p 1mV 5093001p 0mV 5404000p 1mV 5404001p 0mV 5407000p 1mV 5407001p 0mV 5413000p 1mV 5413001p 0mV 5415000p 1mV 5415001p 0mV 5417000p 1mV 5417001p 0mV 5447000p 1mV 5447001p 0mV 5465000p 1mV 5465001p 0mV 5466000p 1mV 5466001p 0mV 5471000p 1mV 5471001p 0mV 5477000p 1mV 5477001p 0mV 5488000p 1mV 5488001p 0mV 5501000p 1mV 5501001p 0mV 5505000p 1mV 5505001p 0mV 5511000p 1mV 5511001p 0mV 5517000p 1mV 5517001p 0mV 5525000p 1mV 5525001p 0mV 5541000p 1mV 5541001p 0mV 5565000p 1mV 5565001p 0mV 5602000p 1mV 5602001p 0mV 5618000p 1mV 5618001p 0mV 5625000p 1mV 5625001p 0mV 5626000p 1mV 5626001p 0mV 5641000p 1mV 5641001p 0mV 5646000p 1mV 5646001p 0mV 5654000p 1mV 5654001p 0mV 5656000p 1mV 5656001p 0mV 5665000p 1mV 5665001p 0mV 5668000p 1mV 5668001p 0mV 5671000p 1mV 5671001p 0mV 5673000p 1mV 5673001p 0mV 5676000p 1mV 5676001p 0mV 5687000p 1mV 5687001p 0mV 5716000p 1mV 5716001p 0mV 5717000p 1mV 5717001p 0mV 5721000p 1mV 5721001p 0mV 5749000p 1mV 5749001p 0mV 5752000p 1mV 5752001p 0mV 5798000p 1mV 5798001p 0mV 5799000p 1mV 5799001p 0mV 5800000p 1mV 5800001p 0mV 5813000p 1mV 5813001p 0mV 5817000p 1mV 5817001p 0mV 5820000p 1mV 5820001p 0mV 5829000p 1mV 5829001p 0mV 5835000p 1mV 5835001p 0mV 5836000p 1mV 5836001p 0mV 5842000p 1mV 5842001p 0mV 5896000p 1mV 5896001p 0mV 5898000p 1mV 5898001p 0mV 5899000p 1mV 5899001p 0mV 6015000p 1mV 6015001p 0mV 6020000p 1mV 6020001p 0mV 6027000p 1mV 6027001p 0mV 6054000p 1mV 6054001p 0mV 6056000p 1mV 6056001p 0mV 6060000p 1mV 6060001p 0mV 6074000p 1mV 6074001p 0mV 6077000p 1mV 6077001p 0mV 6090000p 1mV 6090001p 0mV 6202000p 1mV 6202001p 0mV 6215000p 1mV 6215001p 0mV 6221000p 1mV 6221001p 0mV 6231000p 1mV 6231001p 0mV 6237000p 1mV 6237001p 0mV 6246000p 1mV 6246001p 0mV 6248000p 1mV 6248001p 0mV 6253000p 1mV 6253001p 0mV 6262000p 1mV 6262001p 0mV 6267000p 1mV 6267001p 0mV 6268000p 1mV 6268001p 0mV 6289000p 1mV 6289001p 0mV 6297000p 1mV 6297001p 0mV 6306000p 1mV 6306001p 0mV 6313000p 1mV 6313001p 0mV 6321000p 1mV 6321001p 0mV 6324000p 1mV 6324001p 0mV 6335000p 1mV 6335001p 0mV 6344000p 1mV 6344001p 0mV 6352000p 1mV 6352001p 0mV 6359000p 1mV 6359001p 0mV 6362000p 1mV 6362001p 0mV 6367000p 1mV 6367001p 0mV 6372000p 1mV 6372001p 0mV 6376000p 1mV 6376001p 0mV 6381000p 1mV 6381001p 0mV 6383000p 1mV 6383001p 0mV 6385000p 1mV 6385001p 0mV 6399000p 1mV 6399001p 0mV 6404000p 1mV 6404001p 0mV 6405000p 1mV 6405001p 0mV 6408000p 1mV 6408001p 0mV 6409000p 1mV 6409001p 0mV 6411000p 1mV 6411001p 0mV 6416000p 1mV 6416001p 0mV 6422000p 1mV 6422001p 0mV 6428000p 1mV 6428001p 0mV 6437000p 1mV 6437001p 0mV 6474000p 1mV 6474001p 0mV 6484000p 1mV 6484001p 0mV 6492000p 1mV 6492001p 0mV 6495000p 1mV 6495001p 0mV 6498000p 1mV 6498001p 0mV 6505000p 1mV 6505001p 0mV 6509000p 1mV 6509001p 0mV 6510000p 1mV 6510001p 0mV 6528000p 1mV 6528001p 0mV 6532000p 1mV 6532001p 0mV 6548000p 1mV 6548001p 0mV 6554000p 1mV 6554001p 0mV 6564000p 1mV 6564001p 0mV 6589000p 1mV 6589001p 0mV 6610000p 1mV 6610001p 0mV 6623000p 1mV 6623001p 0mV 6626000p 1mV 6626001p 0mV 6634000p 1mV 6634001p 0mV 6637000p 1mV 6637001p 0mV 6641000p 1mV 6641001p 0mV 6667000p 1mV 6667001p 0mV 6691000p 1mV 6691001p 0mV 6693000p 1mV 6693001p 0mV 6695000p 1mV 6695001p 0mV 6697000p 1mV 6697001p 0mV 6706000p 1mV 6706001p 0mV 6707000p 1mV 6707001p 0mV 6711000p 1mV 6711001p 0mV 6726000p 1mV 6726001p 0mV 6729000p 1mV 6729001p 0mV 6732000p 1mV 6732001p 0mV 6735000p 1mV 6735001p 0mV 6742000p 1mV 6742001p 0mV 6769000p 1mV 6769001p 0mV 6797000p 1mV 6797001p 0mV 6905000p 1mV 6905001p 0mV 6908000p 1mV 6908001p 0mV 6910000p 1mV 6910001p 0mV 6925000p 1mV 6925001p 0mV 6928000p 1mV 6928001p 0mV 6931000p 1mV 6931001p 0mV 6944000p 1mV 6944001p 0mV 6948000p 1mV 6948001p 0mV 6949000p 1mV 6949001p 0mV 6951000p 1mV 6951001p 0mV 6966000p 1mV 6966001p 0mV 6987000p 1mV 6987001p 0mV 6993000p 1mV 6993001p 0mV 6994000p 1mV 6994001p 0mV 6998000p 1mV 6998001p 0mV 7002000p 1mV 7002001p 0mV 7011000p 1mV 7011001p 0mV 7018000p 1mV 7018001p 0mV 7023000p 1mV 7023001p 0mV 7036000p 1mV 7036001p 0mV 7039000p 1mV 7039001p 0mV 7052000p 1mV 7052001p 0mV 7061000p 1mV 7061001p 0mV 7079000p 1mV 7079001p 0mV 7085000p 1mV 7085001p 0mV 7090000p 1mV 7090001p 0mV 7094000p 1mV 7094001p 0mV 7114000p 1mV 7114001p 0mV 7130000p 1mV 7130001p 0mV 7136000p 1mV 7136001p 0mV 7159000p 1mV 7159001p 0mV 7165000p 1mV 7165001p 0mV 7172000p 1mV 7172001p 0mV 7174000p 1mV 7174001p 0mV 7175000p 1mV 7175001p 0mV 7180000p 1mV 7180001p 0mV 7184000p 1mV 7184001p 0mV 7194000p 1mV 7194001p 0mV 7196000p 1mV 7196001p 0mV 7201000p 1mV 7201001p 0mV 7216000p 1mV 7216001p 0mV 7222000p 1mV 7222001p 0mV 7226000p 1mV 7226001p 0mV 7247000p 1mV 7247001p 0mV 7248000p 1mV 7248001p 0mV 7251000p 1mV 7251001p 0mV 7260000p 1mV 7260001p 0mV 7272000p 1mV 7272001p 0mV 7299000p 1mV 7299001p 0mV 7301000p 1mV 7301001p 0mV 7305000p 1mV 7305001p 0mV 7306000p 1mV 7306001p 0mV 7308000p 1mV 7308001p 0mV 7319000p 1mV 7319001p 0mV 7321000p 1mV 7321001p 0mV 7322000p 1mV 7322001p 0mV 7324000p 1mV 7324001p 0mV 7349000p 1mV 7349001p 0mV 7362000p 1mV 7362001p 0mV 7365000p 1mV 7365001p 0mV 7375000p 1mV 7375001p 0mV 7380000p 1mV 7380001p 0mV 7416000p 1mV 7416001p 0mV 7418000p 1mV 7418001p 0mV 7434000p 1mV 7434001p 0mV 7438000p 1mV 7438001p 0mV 7461000p 1mV 7461001p 0mV 7485000p 1mV 7485001p 0mV 7491000p 1mV 7491001p 0mV 7496000p 1mV 7496001p 0mV 7516000p 1mV 7516001p 0mV 7528000p 1mV 7528001p 0mV 7544000p 1mV 7544001p 0mV 7548000p 1mV 7548001p 0mV 7553000p 1mV 7553001p 0mV 7558000p 1mV 7558001p 0mV 7573000p 1mV 7573001p 0mV 7584000p 1mV 7584001p 0mV 7587000p 1mV 7587001p 0mV 7588000p 1mV 7588001p 0mV 7598000p 1mV 7598001p 0mV 7599000p 1mV 7599001p 0mV 7602000p 1mV 7602001p 0mV 7603000p 1mV 7603001p 0mV 7607000p 1mV 7607001p 0mV 7634000p 1mV 7634001p 0mV 7640000p 1mV 7640001p 0mV 7649000p 1mV 7649001p 0mV 7660000p 1mV 7660001p 0mV 7685000p 1mV 7685001p 0mV 7688000p 1mV 7688001p 0mV 7696000p 1mV 7696001p 0mV 7712000p 1mV 7712001p 0mV 7755000p 1mV 7755001p 0mV 7765000p 1mV 7765001p 0mV 7785000p 1mV 7785001p 0mV 7812000p 1mV 7812001p 0mV 7814000p 1mV 7814001p 0mV 7827000p 1mV 7827001p 0mV 7842000p 1mV 7842001p 0mV 7864000p 1mV 7864001p 0mV 7871000p 1mV 7871001p 0mV 7886000p 1mV 7886001p 0mV 7903000p 1mV 7903001p 0mV 7908000p 1mV 7908001p 0mV 7909000p 1mV 7909001p 0mV 7918000p 1mV 7918001p 0mV 7922000p 1mV 7922001p 0mV 7927000p 1mV 7927001p 0mV 7930000p 1mV 7930001p 0mV 7951000p 1mV 7951001p 0mV 7968000p 1mV 7968001p 0mV 7985000p 1mV 7985001p 0mV 7988000p 1mV 7988001p 0mV 7990000p 1mV 7990001p 0mV 8012000p 1mV 8012001p 0mV 8014000p 1mV 8014001p 0mV 8040000p 1mV 8040001p 0mV 8043000p 1mV 8043001p 0mV 8050000p 1mV 8050001p 0mV 8057000p 1mV 8057001p 0mV 8067000p 1mV 8067001p 0mV 8084000p 1mV 8084001p 0mV 8086000p 1mV 8086001p 0mV 8098000p 1mV 8098001p 0mV 8129000p 1mV 8129001p 0mV 8137000p 1mV 8137001p 0mV 8148000p 1mV 8148001p 0mV 8155000p 1mV 8155001p 0mV 8158000p 1mV 8158001p 0mV 8164000p 1mV 8164001p 0mV 8167000p 1mV 8167001p 0mV 8176000p 1mV 8176001p 0mV 8187000p 1mV 8187001p 0mV 8189000p 1mV 8189001p 0mV 8203000p 1mV 8203001p 0mV 8206000p 1mV 8206001p 0mV 8208000p 1mV 8208001p 0mV 8214000p 1mV 8214001p 0mV 8219000p 1mV 8219001p 0mV 8227000p 1mV 8227001p 0mV 8271000p 1mV 8271001p 0mV 8301000p 1mV 8301001p 0mV 8307000p 1mV 8307001p 0mV 8309000p 1mV 8309001p 0mV 8319000p 1mV 8319001p 0mV 8321000p 1mV 8321001p 0mV 8323000p 1mV 8323001p 0mV 8337000p 1mV 8337001p 0mV 8338000p 1mV 8338001p 0mV 8341000p 1mV 8341001p 0mV 8342000p 1mV 8342001p 0mV 8347000p 1mV 8347001p 0mV 8362000p 1mV 8362001p 0mV 8372000p 1mV 8372001p 0mV 8381000p 1mV 8381001p 0mV 8416000p 1mV 8416001p 0mV 8445000p 1mV 8445001p 0mV 8457000p 1mV 8457001p 0mV 8473000p 1mV 8473001p 0mV 8479000p 1mV 8479001p 0mV 8493000p 1mV 8493001p 0mV 8503000p 1mV 8503001p 0mV 8505000p 1mV 8505001p 0mV 8523000p 1mV 8523001p 0mV 8536000p 1mV 8536001p 0mV 8537000p 1mV 8537001p 0mV 8548000p 1mV 8548001p 0mV 8561000p 1mV 8561001p 0mV 8564000p 1mV 8564001p 0mV 8566000p 1mV 8566001p 0mV 8587000p 1mV 8587001p 0mV 8598000p 1mV 8598001p 0mV 8605000p 1mV 8605001p 0mV 8613000p 1mV 8613001p 0mV 8624000p 1mV 8624001p 0mV 8627000p 1mV 8627001p 0mV 8628000p 1mV 8628001p 0mV 8630000p 1mV 8630001p 0mV 8641000p 1mV 8641001p 0mV 8650000p 1mV 8650001p 0mV 8655000p 1mV 8655001p 0mV 8659000p 1mV 8659001p 0mV 8664000p 1mV 8664001p 0mV 8668000p 1mV 8668001p 0mV 8671000p 1mV 8671001p 0mV 8683000p 1mV 8683001p 0mV 8684000p 1mV 8684001p 0mV 8701000p 1mV 8701001p 0mV 8711000p 1mV 8711001p 0mV 8744000p 1mV 8744001p 0mV 8754000p 1mV 8754001p 0mV 8760000p 1mV 8760001p 0mV 8762000p 1mV 8762001p 0mV 8791000p 1mV 8791001p 0mV 8793000p 1mV 8793001p 0mV 8908000p 1mV 8908001p 0mV 8918000p 1mV 8918001p 0mV 8923000p 1mV 8923001p 0mV 8951000p 1mV 8951001p 0mV 8953000p 1mV 8953001p 0mV 8973000p 1mV 8973001p 0mV 8975000p 1mV 8975001p 0mV 8982000p 1mV 8982001p 0mV 8999000p 1mV 8999001p 0mV 9008000p 1mV 9008001p 0mV 9009000p 1mV 9009001p 0mV 9016000p 1mV 9016001p 0mV 9020000p 1mV 9020001p 0mV 9028000p 1mV 9028001p 0mV 9038000p 1mV 9038001p 0mV 9044000p 1mV 9044001p 0mV 9068000p 1mV 9068001p 0mV 9074000p 1mV 9074001p 0mV 9076000p 1mV 9076001p 0mV 9092000p 1mV 9092001p 0mV 9093000p 1mV 9093001p 0mV 9098000p 1mV 9098001p 0mV 9112000p 1mV 9112001p 0mV 9116000p 1mV 9116001p 0mV 9117000p 1mV 9117001p 0mV 9118000p 1mV 9118001p 0mV 9156000p 1mV 9156001p 0mV 9163000p 1mV 9163001p 0mV 9164000p 1mV 9164001p 0mV 9180000p 1mV 9180001p 0mV 9191000p 1mV 9191001p 0mV 9204000p 1mV 9204001p 0mV 9205000p 1mV 9205001p 0mV 9217000p 1mV 9217001p 0mV 9218000p 1mV 9218001p 0mV 9220000p 1mV 9220001p 0mV 9251000p 1mV 9251001p 0mV 9260000p 1mV 9260001p 0mV 9274000p 1mV 9274001p 0mV 9289000p 1mV 9289001p 0mV 9304000p 1mV 9304001p 0mV 9319000p 1mV 9319001p 0mV 9327000p 1mV 9327001p 0mV 9334000p 1mV 9334001p 0mV 9365000p 1mV 9365001p 0mV 9407000p 1mV 9407001p 0mV 9410000p 1mV 9410001p 0mV 9421000p 1mV 9421001p 0mV 9429000p 1mV 9429001p 0mV 9431000p 1mV 9431001p 0mV 9441000p 1mV 9441001p 0mV 9457000p 1mV 9457001p 0mV 9484000p 1mV 9484001p 0mV 9489000p 1mV 9489001p 0mV 9490000p 1mV 9490001p 0mV 9495000p 1mV 9495001p 0mV 9507000p 1mV 9507001p 0mV 9518000p 1mV 9518001p 0mV 9525000p 1mV 9525001p 0mV 9530000p 1mV 9530001p 0mV 9536000p 1mV 9536001p 0mV 9546000p 1mV 9546001p 0mV 9553000p 1mV 9553001p 0mV 9563000p 1mV 9563001p 0mV 9564000p 1mV 9564001p 0mV)
.ENDS conductors__anyBias-Lk_0_704



XVI1 28 285 conductors__anyBias-Lk_0_701
XREF1 B1 285 gnd newJTL__phaseReference
RR1  28 285 100

XVI2  37 385 conductors__anyBias-Lk_0_702
XREF2 B2 385 gnd newJTL__phaseReference
RR2  37 385 100

XVI3  64 485 conductors__anyBias-Lk_0_703
XREF3 B3 485 gnd newJTL__phaseReference
RR3  64 485 100

XVI4  73  585 conductors__anyBias-Lk_0_704
XREF4 B4 585 gnd newJTL__phaseReference
RR4 73  585  100






****TOP LEVEL CELL: aNewTestLibrary:testJTL{sch}


XJ1 1 junctionsBypassGround__gbj1p0
Xbias1 1 conductors__anyBias-Lk_0
XLL1 1 2 inductors__fixedInd1p5
XJ2 2 junctionsBypassGround__gbj1p0
Xbias2 2 conductors__anyBias-Lk_0
XLL2 2 3 inductors__fixedInd1p5
XJ3 3 junctionsBypassGround__gbj1p0
Xbias3 3 conductors__anyBias-Lk_0
XLL3 3 4 inductors__fixedInd1p5
XJ4 4 junctionsBypassGround__gbj1p0
Xbias4 4 conductors__anyBias-Lk_0
XLL4 4 5 inductors__fixedInd1p5
XJ5 5 junctionsBypassGround__gbj1p0
Xbias5 5 conductors__anyBias-Lk_0
XLL5 5 6 inductors__fixedInd1p5
XJ6 6 junctionsBypassGround__gbj1p0
Xbias6 6 conductors__anyBias-Lk_0
XLL6 6 7 inductors__fixedInd1p5
XJ7 7 junctionsBypassGround__gbj1p0
Xbias7 7 conductors__anyBias-Lk_0
XLL7 7 8 inductors__fixedInd1p5
XJ8 8 junctionsBypassGround__gbj1p0
Xbias8 8 conductors__anyBias-Lk_0
XLL8 8 9 inductors__fixedInd1p5
XJ9 9 junctionsBypassGround__gbj1p0
Xbias9 9 conductors__anyBias-Lk_0

XLL100 1 11 inductors__fixedInd1p5
XLL200 2 12 inductors__fixedInd1p5
XLL300 3 13 inductors__fixedInd1p5
XLL400 4 14 inductors__fixedInd1p5
XLL500 5 15 inductors__fixedInd1p5
XLL600 6 16 inductors__fixedInd1p5
XLL700 7 17 inductors__fixedInd1p5
XLL800 8 18 inductors__fixedInd1p5
XLL900 9 19 inductors__fixedInd1p5


XJ10 11 junctionsBypassGround__gbj1p0
Xbias10 11 conductors__anyBias-Lk_0
XLL10 11 12 inductors__fixedInd1p5
XJ11 12 junctionsBypassGround__gbj1p0
Xbias11 12 conductors__anyBias-Lk_0
XLL11 12 13 inductors__fixedInd1p5
XJ12 13 junctionsBypassGround__gbj1p0
Xbias12 13 conductors__anyBias-Lk_0
XLL12 13 14 inductors__fixedInd1p5
XJ13 14 junctionsBypassGround__gbj1p0
Xbias13 14 conductors__anyBias-Lk_0
XLL13 14 15 inductors__fixedInd1p5
XJ14 15 junctionsBypassGround__gbj1p0
Xbias14 15 conductors__anyBias-Lk_0
XLL14 15 16 inductors__fixedInd1p5
XJ15 16 junctionsBypassGround__gbj1p0
Xbias15 16 conductors__anyBias-Lk_0
XLL15 16 17 inductors__fixedInd1p5
XJ16 17 junctionsBypassGround__gbj1p0
Xbias16 17 conductors__anyBias-Lk_0
XLL16 17 18 inductors__fixedInd1p5
XJ17 18 junctionsBypassGround__gbj1p0
Xbias17 18 conductors__anyBias-Lk_0
XLL17 17 18 inductors__fixedInd1p5
XJ18 19 junctionsBypassGround__gbj1p0
Xbias18 19 conductors__anyBias-Lk_0

XLL110  11 21 inductors__fixedInd1p5
XLL210  12 22 inductors__fixedInd1p5
XLL310  13 23 inductors__fixedInd1p5
XLL410  14 24 inductors__fixedInd1p5
XLL510  15 25 inductors__fixedInd1p5
XLL610  16 26 inductors__fixedInd1p5
XLL710  17 27 inductors__fixedInd1p5
XLL810  18 28 inductors__fixedInd1p5
XLL910  19 29 inductors__fixedInd1p5

XJ19 21 junctionsBypassGround__gbj1p0
XLL19 21 22 inductors__fixedInd1p5
Xbias19 21 conductors__anyBias-Lk_0
XJ20 22 junctionsBypassGround__gbj1p0
Xbias20 22 conductors__anyBias-Lk_0
XLL20 22 23 inductors__fixedInd1p5
XJ21 23 junctionsBypassGround__gbj1p0
XLL21 23 24 inductors__fixedInd1p5
Xbias21 23 conductors__anyBias-Lk_0
XJ22 24 junctionsBypassGround__gbj1p0
Xbias22 24 conductors__anyBias-Lk_0
XLL22 24 25 inductors__fixedInd1p5
XJ23 25 junctionsBypassGround__gbj1p0
Xbias23 25 conductors__anyBias-Lk_0
XLL23 25 26 inductors__fixedInd1p5
XJ24 26 junctionsBypassGround__gbj1p0
Xbias24 26 conductors__anyBias-Lk_0
XLL24 26 27 inductors__fixedInd1p5
XJ25 27 junctionsBypassGround__gbj1p0
Xbias25 27 conductors__anyBias-Lk_0
XLL25 27 28 inductors__fixedInd1p5
XJ26 28 junctionsBypassGround__gbj1p0
Xbias26 28 conductors__anyBias-Lk_0
XLL26 28 29 inductors__fixedInd1p5
XJ27 29 junctionsBypassGround__gbj1p0
Xbias27 29 conductors__anyBias-Lk_0

XLL120   21 31 inductors__fixedInd1p5
XLL220   22 32 inductors__fixedInd1p5
XLL320   23 33 inductors__fixedInd1p5
XLL420   24 34 inductors__fixedInd1p5
XLL520   25 35 inductors__fixedInd1p5
XLL620   26 36 inductors__fixedInd1p5
XLL720   27 37 inductors__fixedInd1p5
XLL820   28 38 inductors__fixedInd1p5
XLL920   29 39 inductors__fixedInd1p5


XJ28 31 junctionsBypassGround__gbj1p0
XLL28 31 32 inductors__fixedInd1p5
Xbias28 31 conductors__anyBias-Lk_0
XJ29 32 junctionsBypassGround__gbj1p0
Xbias29 32 conductors__anyBias-Lk_0
XLL29 32 33 inductors__fixedInd1p5
XJ30 33 junctionsBypassGround__gbj1p0
XLL30 33 34 inductors__fixedInd1p5
Xbias30 33 conductors__anyBias-Lk_0
XJ31 34 junctionsBypassGround__gbj1p0
Xbias31 34 conductors__anyBias-Lk_0
XLL31 34 35 inductors__fixedInd1p5
XJ32 35 junctionsBypassGround__gbj1p0
Xbias32 35 conductors__anyBias-Lk_0
XLL32 35 36 inductors__fixedInd1p5
XJ33 36 junctionsBypassGround__gbj1p0
Xbias33 36 conductors__anyBias-Lk_0
XLL33 36 37 inductors__fixedInd1p5
XJ34 37 junctionsBypassGround__gbj1p0
Xbias34 37 conductors__anyBias-Lk_0
XLL34 37 38 inductors__fixedInd1p5
XJ35 38 junctionsBypassGround__gbj1p0
Xbias35 38 conductors__anyBias-Lk_0
XLL35 38 39 inductors__fixedInd1p5
XJ36 39 junctionsBypassGround__gbj1p0
Xbias36 39 conductors__anyBias-Lk_0


XLL130  31 41 inductors__fixedInd1p5
XLL230  32 42 inductors__fixedInd1p5
XLL330  33 43 inductors__fixedInd1p5
XLL430  34 44 inductors__fixedInd1p5
XLL530  35 45 inductors__fixedInd1p5
XLL630  36 46 inductors__fixedInd1p5
XLL730  37 47 inductors__fixedInd1p5
XLL830  38 48 inductors__fixedInd1p5
XLL930  39 49 inductors__fixedInd1p5



XJ37 41 junctionsBypassGround__gbj1p0
Xbias37 41 conductors__anyBias-Lk_0
XLL37 41 42 inductors__fixedInd1p5
XJ38 42 junctionsBypassGround__gbj1p0
Xbias38 42 conductors__anyBias-Lk_0
XLL38 42 43 inductors__fixedInd1p5
XJ39 43 junctionsBypassGround__gbj1p0
Xbias39 43 conductors__anyBias-Lk_0
XLL39 43 44 inductors__fixedInd1p5
XJ40 44 junctionsBypassGround__gbj1p0
Xbias40 44 conductors__anyBias-Lk_0
XLL40 44 45 inductors__fixedInd1p5
XJ41 45 junctionsBypassGround__gbj1p0
Xbias41 45 conductors__anyBias-Lk_0
XLL41 45 46 inductors__fixedInd1p5
XJ42 46 junctionsBypassGround__gbj1p0
Xbias42 46 conductors__anyBias-Lk_0
XLL42 46 47 inductors__fixedInd1p5
XJ43 47 junctionsBypassGround__gbj1p0
Xbias43 47 conductors__anyBias-Lk_0
XLL43 47 48 inductors__fixedInd1p5
XJ44 48 junctionsBypassGround__gbj1p0
Xbias44 48 conductors__anyBias-Lk_0
XLL44 48 49 inductors__fixedInd1p5
XJ45 49 junctionsBypassGround__gbj1p0
Xbias45 49 conductors__anyBias-Lk_0


XLL140  41 51 inductors__fixedInd1p5
XLL240  42 52 inductors__fixedInd1p5
XLL340  43 53 inductors__fixedInd1p5
XLL440  44 54 inductors__fixedInd1p5
XLL540  45 55 inductors__fixedInd1p5
XLL640  46 56 inductors__fixedInd1p5
XLL740  47 57 inductors__fixedInd1p5
XLL840  48 58 inductors__fixedInd1p5
XLL940  49 59 inductors__fixedInd1p5

XJ46 51 junctionsBypassGround__gbj1p0
Xbias46 51 conductors__anyBias-Lk_0
XLL46 51 52 inductors__fixedInd1p5
XJ47 52 junctionsBypassGround__gbj1p0
Xbias47 52 conductors__anyBias-Lk_0
XLL47 52 53 inductors__fixedInd1p5
XJ48 53 junctionsBypassGround__gbj1p0
Xbias48 53 conductors__anyBias-Lk_0
XLL48 53 54 inductors__fixedInd1p5
XJ49 54 junctionsBypassGround__gbj1p0
Xbias49 54 conductors__anyBias-Lk_0
XLL49 54 55 inductors__fixedInd1p5
XJ50 55 junctionsBypassGround__gbj1p0
Xbias50 55 conductors__anyBias-Lk_0
XLL50 55 56 inductors__fixedInd1p5
XJ51 56 junctionsBypassGround__gbj1p0
Xbias51 56 conductors__anyBias-Lk_0
XLL51 56 57 inductors__fixedInd1p5
XJ52 57 junctionsBypassGround__gbj1p0
Xbias52 57 conductors__anyBias-Lk_0
XLL52 57 58 inductors__fixedInd1p5
XJ53 58 junctionsBypassGround__gbj1p0
Xbias53 58 conductors__anyBias-Lk_0
XLL53 58 59 inductors__fixedInd1p5
XJ54 59 junctionsBypassGround__gbj1p0
Xbias54 59 conductors__anyBias-Lk_0

XLL150  51 61 inductors__fixedInd1p5
XLL250  52 62 inductors__fixedInd1p5
XLL350  53 63 inductors__fixedInd1p5
XLL450  54 64 inductors__fixedInd1p5
XLL550  55 65 inductors__fixedInd1p5
XLL650  56 66 inductors__fixedInd1p5
XLL750  57 67 inductors__fixedInd1p5
XLL850  58 68 inductors__fixedInd1p5
XLL950  59 69 inductors__fixedInd1p5

XJ55 61 junctionsBypassGround__gbj1p0
Xbias55 61 conductors__anyBias-Lk_0
XLL55 61 62 inductors__fixedInd1p5
XJ56 62 junctionsBypassGround__gbj1p0
Xbias56 62 conductors__anyBias-Lk_0
XLL56 62 63 inductors__fixedInd1p5
XJ57 63 junctionsBypassGround__gbj1p0
Xbias57 63 conductors__anyBias-Lk_0
XLL57 63 64 inductors__fixedInd1p5
XJ58 64 junctionsBypassGround__gbj1p0
Xbias58 64 conductors__anyBias-Lk_0
XLL58 64 65 inductors__fixedInd1p5
XJ59 65 junctionsBypassGround__gbj1p0
Xbias59 65 conductors__anyBias-Lk_0
XLL59 65 66 inductors__fixedInd1p5
XJ60 66 junctionsBypassGround__gbj1p0
Xbias60 66 conductors__anyBias-Lk_0
XLL60 66 67 inductors__fixedInd1p5
XJ61 67 junctionsBypassGround__gbj1p0
Xbias61 67 conductors__anyBias-Lk_0
XLL61 67 68 inductors__fixedInd1p5
XJ62 68 junctionsBypassGround__gbj1p0
Xbias62 68 conductors__anyBias-Lk_0
XLL62 68 69 inductors__fixedInd1p5
XJ63 69 junctionsBypassGround__gbj1p0
Xbias63 69 conductors__anyBias-Lk_0


XLL160  61 71 inductors__fixedInd1p5
XLL260  62 72 inductors__fixedInd1p5
XLL360  63 73 inductors__fixedInd1p5
XLL460  64 74 inductors__fixedInd1p5
XLL560  65 75 inductors__fixedInd1p5
XLL660  66 76 inductors__fixedInd1p5
XLL760  67 77 inductors__fixedInd1p5
XLL860  68 78 inductors__fixedInd1p5
XLL960  69 79 inductors__fixedInd1p5


XJ64 71 junctionsBypassGround__gbj1p0
Xbias64 71 conductors__anyBias-Lk_0
XLL64 71 72 inductors__fixedInd1p5
XJ65 72 junctionsBypassGround__gbj1p0
Xbias65 72 conductors__anyBias-Lk_0
XLL65 72 73 inductors__fixedInd1p5
XJ66 73 junctionsBypassGround__gbj1p0
Xbias66 73 conductors__anyBias-Lk_0
XLL66 73 74 inductors__fixedInd1p5
XJ67 74 junctionsBypassGround__gbj1p0
Xbias67 74 conductors__anyBias-Lk_0
XLL67 74 75 inductors__fixedInd1p5
XJ68 75 junctionsBypassGround__gbj1p0
Xbias68 75 conductors__anyBias-Lk_0
XLL68 75 76 inductors__fixedInd1p5
XJ69 76 junctionsBypassGround__gbj1p0
Xbias69 76 conductors__anyBias-Lk_0
XLL69 76 77 inductors__fixedInd1p5
XJ70 77 junctionsBypassGround__gbj1p0
Xbias70 77 conductors__anyBias-Lk_0
XLL70 77 78 inductors__fixedInd1p5
XJ71 78 junctionsBypassGround__gbj1p0
Xbias71 78 conductors__anyBias-Lk_0
XLL71 78 79 inductors__fixedInd1p5
XJ72 79 junctionsBypassGround__gbj1p0
Xbias72 79 conductors__anyBias-Lk_0


XLL170  71 81 inductors__fixedInd1p5
XLL270  72 82 inductors__fixedInd1p5
XLL370  73 83 inductors__fixedInd1p5
XLL470  74 84 inductors__fixedInd1p5
XLL570  75 85 inductors__fixedInd1p5
XLL670  76 86 inductors__fixedInd1p5
XLL770  77 87 inductors__fixedInd1p5
XLL870  78 88 inductors__fixedInd1p5
XLL970  79 89 inductors__fixedInd1p5


XJ73 81 junctionsBypassGround__gbj1p0
Xbias73 81 conductors__anyBias-Lk_0
XLL73 81 82 inductors__fixedInd1p5
XJ74 82 junctionsBypassGround__gbj1p0
Xbias74 82 conductors__anyBias-Lk_0
XLL74 82 83 inductors__fixedInd1p5
XJ75 83 junctionsBypassGround__gbj1p0
Xbias75 83 conductors__anyBias-Lk_0
XLL75 83 84 inductors__fixedInd1p5
XJ76 84 junctionsBypassGround__gbj1p0
Xbias76 84 conductors__anyBias-Lk_0
XLL76 84 85 inductors__fixedInd1p5
XJ77 85 junctionsBypassGround__gbj1p0
Xbias77 85 conductors__anyBias-Lk_0
XLL77 85 86 inductors__fixedInd1p5
XJ78 86 junctionsBypassGround__gbj1p0
Xbias78 86 conductors__anyBias-Lk_0
XLL78 86 87 inductors__fixedInd1p5
XJ79 87 junctionsBypassGround__gbj1p0
Xbias79 87 conductors__anyBias-Lk_0
XLL79 87 88 inductors__fixedInd1p5
XJ80 89 junctionsBypassGround__gbj1p0
Xbias80 89 conductors__anyBias-Lk_0
XLL80 89 90 inductors__fixedInd1p5
XJ81 91 junctionsBypassGround__gbj1p0
Xbias81 91 conductors__anyBias-Lk_0

.END
