*** SPICE deck for cell testJTLplain{sch} from library aNewTestLibrary
*** Created on Sat Jan 09, 2021 14:13:09
*** Last revised on Mon Aug 26, 2024 11:38:12
*** Written on Mon Aug 26, 2024 11:55:08 by Electric VLSI Design System, version 9.08e
*** Layout tech: josephson, foundry NONE
*** UC SPICE *** , MIN_RESIST 0.0, MIN_CAPAC 0.0FF
* Model cards copied from file: /Users/ivans/years/2020-2024/2024/2024-ivan/electric-2024/theBest1aug24/aTests/testJTLplain.txt
*** These are the print statement for testJTLplain
*** ies 26 August 2024
*** josim -o Aoutput.csv testJTLplain.cir 



.tran 0.1p 100p 0 0.1p


.print DEVV BJi|xJ36
.print DEVV BJi|xJ37
.print DEVV BJi|xJ64
.print DEVV BJi|xJ73




* End of Model cards copied from file: /Users/ivans/years/2020-2024/2024/2024-ivan/electric-2024/theBest1jul24/aTests/testJTL.txt
.model jmitll jj(rtype=1, vg=.002V, cap=0.07pF, r0=160, rN=16, icrit=0.0001A)


.SUBCKT junctionsBypassGround__gbj1p0 D 
BJi D gnd jmitll area=1.25
RRi D gnd 5.36
.ENDS junctionsBypassGround__gbj1p0


*** SUBCIRCUIT inductors__fixedInd1p5 FROM CELL inductors:fixedInd3p0{sch}
.SUBCKT inductors__fixedInd1p5 A B
LLi A B 7.891E-12
.ENDS inductors__fixedInd1p5


*** SUBCIRCUIT conductors__anyBias-Lk_0 FROM CELL conductors:anyBias{sch}
.SUBCKT conductors__anyBias-Lk_0  D
RR1 NN D 29.42
VrampSppl@0 NN gnd pwl (0 0 1p 0.0026V)
.ENDS conductors__anyBias-Lk_0_707



****.SUBCKT conductors__anyBias-Lk_0 D
****RR1 NN D 8
****VrampSppl@0 NN gnd pwl (0 0 1p 3.86V)
***.ENDS conductors__anyBias-Lk_0

*** SUBCIRCUIT junctions__jb2p0 FROM CELL junctions:jb2p0{sch}
.SUBCKT junctions__jb2p0 D S
BJi S D jmitll area=2.5
RRi S D 2.68
.ENDS junctions__jb2p0

*** SUBCIRCUIT junctions__jb200p0 FROM CELL junctions:jb200p0{sch}
.SUBCKT junctions__jb200p0 D S
BJi S D jmitll area=250.0
RRi S D 0.0268
.ENDS junctions__jb200p0

*** SUBCIRCUIT conductors__anyBias-Lk_1_414 FROM CELL conductors:anyBias{sch}
.SUBCKT conductors__anyBias-Lk_1_414 D
RR1 NN D 14.71
VrampSppl@0 NN gnd pwl (0 0 1p 0.0026V)
.ENDS conductors__anyBias-Lk_1_414

*** SUBCIRCUIT conductors__bias1p4 FROM CELL conductors:bias1p4{sch}
.SUBCKT conductors__bias1p4 D
Xnormaliz@0 D conductors__anyBias-Lk_1_414
.ENDS conductors__bias1p4

*** SUBCIRCUIT conductors__anyBias-Lk_141_4 FROM CELL conductors:anyBias{sch}
.SUBCKT conductors__anyBias-Lk_141_4 D
RR1 NN D 0.147
VrampSppl@0 NN gnd pwl (0 0 1p 0.0026V)
.ENDS conductors__anyBias-Lk_141_4

*** SUBCIRCUIT conductors__bias1p4x100 FROM CELL conductors:bias1p4x100{sch}
.SUBCKT conductors__bias1p4x100 D
Xnormaliz@0 D conductors__anyBias-Lk_141_4
.ENDS conductors__bias1p4x100

*** SUBCIRCUIT newJTL__phaseReference FROM CELL newJTL:phaseReference{sch}
.SUBCKT newJTL__phaseReference B1 B2 gnd
XJ1 gnd B1 junctions__jb2p0
XJ2 gnd B2 junctions__jb200p0
LM1 net@4 B1 10e-16
LM2 net@3 B2 10e-16
Xbias1p4@0 net@4 conductors__bias1p4
Xbias1p4x@0 net@3 conductors__bias1p4x100
.ENDS newJTL__phaseReference



**cart_pole_input**
.SUBCKT conductors__anyBias-Lk_0_701 bottom out
VrampSppl@0 bottom out pwl (0 0 53.042p 0.553245mV 1007.368p 0.547385mV 1007.631p 0.547385mV 1032.356p 0.550323mV 1045.228p 0.556041mV 1058.556p 0.560958mV 2037.202p 0.553138mV 2056.869p 0.550142mV 2057.657p 0.550142mV 2060.563p 0.549759mV 2094.984p 0.550728mV 2108.134p 0.552483mV 2117.083p 0.554992mV 2126.923p 0.558967mV 2133.567p 0.561505mV 3011.392p 0.551276mV 3020.87p 0.550888mV 3024.101p 0.550888mV 4006.911p 0.550233mV 4010.238p 0.550567mV 4010.649p 0.550567mV 4019.206p 0.550533mV 4019.303p 0.550533mV 4020.943p 0.550133mV 4031.1p 0.548232mV 4038.276p 0.547462mV 4041.034p 0.546325mV 5002.691p 0.553369mV 5020.594p 0.553419mV 5047.768p 0.554227mV 5072.396p 0.551037mV 5111.032p 0.540957mV 6022.417p 0.551098mV 6046.535p 0.550651mV 6059.294p 0.548205mV 6064.527p 0.547164mV 6069.594p 0.545755mV 6083.229p 0.540056mV 7017.643p 0.553323mV 7042.447p 0.551113mV 7051.511p 0.5516mV 7062.419p 0.552074mV 7094.687p 0.557068mV 7129.723p 0.556842mV 8004.237p 0.550534mV 8028.837p 0.552338mV 8050.54p 0.552347mV 8081.527p 0.548688mV 8104.424p 0.541886mV 8115.954p 0.536233mV 9007.123p 0.551225mV 9008.942p 0.551225mV 9026.814p 0.554118mV 9027.223p 0.554118mV 9053.738p 0.55812mV 9061.123p 0.560686mV 10001.474p 0.548939mV 10043.312p 0.538707mV 11057.086p 0.558893mV 11065.573p 0.562009mV 12020.228p 0.554004mV 12041.683p 0.54966mV 12046.602p 0.548935mV 12057.286p 0.548573mV 12058.752p 0.548573mV 12076.955p 0.547806mV 12088.01p 0.547399mV 13045.316p 0.542993mV 13046.642p 0.542993mV 13063.574p 0.540567mV 13081.382p 0.536575mV 14000.139p 0.546113mV 14020.055p 0.54649mV 14021.821p 0.54649mV 14030.804p 0.545941mV 14039.956p 0.545848mV 15031.469p 0.548293mV 15044.659p 0.547114mV 15064.025p 0.545464mV 15075.478p 0.54274mV 15087.162p 0.540056mV 16000.435p 0.552884mV 16012.296p 0.553095mV 16030.639p 0.55353mV 16038.748p 0.552728mV 17031.823p 0.551033mV 17042.498p 0.552093mV 17046.626p 0.552808mV 18052.335p 0.544544mV 18057.381p 0.544514mV 18067.973p 0.54481mV 18072.723p 0.544405mV 19003.008p 0.552928mV 19033.074p 0.549988mV 19034.341p 0.549988mV 19063.306p 0.54559mV 19087.259p 0.540119mV 20019.817p 0.551014mV 20046.995p 0.546428mV 21024.173p 0.549339mV 21026.12p 0.549276mV 21026.489p 0.549276mV 21049.556p 0.548291mV 21056.533p 0.549263mV 21060.436p 0.550297mV 22007.836p 0.554077mV 22028.031p 0.552843mV 22031.752p 0.552534mV 22081.493p 0.5461mV 22116.731p 0.55397mV 22118.004p 0.55397mV 22122.632p 0.555813mV 22147.67p 0.569771mV 22148.893p 0.569771mV 22152.471p 0.572345mV 22153.688p 0.572345mV 23016.269p 0.548965mV 23025.952p 0.549375mV 23041.252p 0.549447mV 23046.334p 0.548741mV 23082.46p 0.541613mV 23096.494p 0.53619mV 23103.282p 0.533646mV 24002.885p 0.54841mV 24025.457p 0.551821mV 24039.768p 0.555757mV 25009.947p 0.548268mV 25028.045p 0.547673mV 25031.108p 0.547343mV 25039.809p 0.547379mV 25045.133p 0.547819mV 25059.849p 0.548992mV 25063.903p 0.549397mV 25068.206p 0.549437mV 25103.31p 0.548289mV 25114.485p 0.546561mV 26000.139p 0.55216mV 26005.459p 0.552106mV 26013.226p 0.552417mV 26022.179p 0.554136mV 26043.789p 0.555384mV 26059.997p 0.555602mV 26078.539p 0.553963mV 26079.396p 0.553963mV 26081.033p 0.553557mV 26091.805p 0.553848mV 27038.009p 0.551694mV 27051.315p 0.556002mV 27063.204p 0.558515mV 27066.188p 0.559959mV 28003.87p 0.551146mV 28015.866p 0.552306mV 28052.094p 0.554626mV 28072.421p 0.562742mV 28073.938p 0.562742mV 28078.067p 0.564958mV 30034.828p 0.54941mV 30063.942p 0.55435mV 30076.045p 0.55629mV 30083.98p 0.556697mV 30100.318p 0.554701mV 30153.714p 0.53739mV 31027.423p 0.548161mV 31124.165p 0.561413mV 32025.143p 0.543779mV 32034.899p 0.543331mV 32038.872p 0.54325mV 32047.129p 0.542724mV 32047.429p 0.542724mV 32054.336p 0.54228mV 33023.594p 0.550992mV 33091.049p 0.547449mV 33107.908p 0.541759mV 33112.322p 0.539858mV 34005.837p 0.554288mV 34007.423p 0.554288mV 34028.976p 0.554303mV 34038.135p 0.553222mV 34066.209p 0.551467mV 34095.826p 0.553399mV 34102.437p 0.554517mV 34133.37p 0.556535mV 34136.225p 0.55658mV 34143.118p 0.556265mV 34146.798p 0.555589mV 34163.907p 0.551404mV 34167.024p 0.549289mV 34194.568p 0.538403mV 34207.335p 0.531757mV 34228.313p 0.521205mV 34261.274p 0.506549mV 34271.086p 0.500515mV 35021.935p 0.548214mV 35022.289p 0.548214mV 35049.774p 0.552594mV 35064.942p 0.555533mV 35088.193p 0.556363mV 35096.92p 0.55607mV 36041.608p 0.546962mV 36055.099p 0.545347mV 36077.808p 0.542677mV 36083.622p 0.542367mV 37011.556p 0.551059mV 37012.909p 0.551059mV 37037.55p 0.549293mV 37043.173p 0.548282mV 37053.853p 0.546626mV 37074.89p 0.541838mV 38017.349p 0.55155mV 38040.47p 0.54797mV 38077.979p 0.544538mV 38081.027p 0.543519mV 39031.22p 0.549651mV 39091.499p 0.555774mV 39158.482p 0.564286mV 39171.229p 0.563023mV 40003.392p 0.551946mV 40016.229p 0.551309mV 40067.595p 0.552193mV 40107.245p 0.555819mV 40131.409p 0.557203mV 40177.102p 0.549962mV 40183.417p 0.5488mV 40215.471p 0.542131mV 40248.445p 0.538422mV 40249.855p 0.538422mV 41020.461p 0.550736mV 41047.327p 0.553302mV 41047.558p 0.553302mV 41069.591p 0.554318mV 41077.588p 0.55336mV 41080.735p 0.552331mV 41108.167p 0.54826mV 41111.575p 0.547218mV 41119.54p 0.546538mV 43033.019p 0.546556mV 43033.024p 0.546556mV 43033.123p 0.546556mV 43040.331p 0.546971mV 43042.821p 0.546971mV 43061.242p 0.549279mV 43068.775p 0.549313mV 43075.22p 0.549753mV 43089.894p 0.550935mV 43098.188p 0.551399mV 43107.126p 0.550418mV 43121.887p 0.5477mV 43137.926p 0.543923mV 43143.356p 0.542915mV 43171.57p 0.532185mV 43183.572p 0.526922mV 44031.713p 0.546297mV 45010.801p 0.551498mV 45010.895p 0.551498mV 46008.214p 0.546274mV 46051.02p 0.542256mV 46057.836p 0.541522mV 46072.798p 0.539313mV 46076.112p 0.538572mV 46098.557p 0.53558mV 47002.05p 0.553095mV 47022.04p 0.553001mV 47023.994p 0.553001mV 47024.201p 0.553001mV 47031.823p 0.553323mV 47103.822p 0.545437mV 47105.924p 0.543962mV 47106.648p 0.543962mV 48049.351p 0.559991mV 49000.774p 0.553413mV 49044.289p 0.555502mV 49049.416p 0.555496mV 49057.852p 0.555855mV 49069.026p 0.556225mV 49088.483p 0.557728mV 49093.255p 0.558843mV 50018.916p 0.550154mV 50029.549p 0.549881mV 50039.587p 0.550341mV 50042.02p 0.550754mV 50048.219p 0.551533mV 50065.247p 0.553195mV 50097.6p 0.55244mV 50099.283p 0.55244mV 50100.348p 0.551406mV 50117.358p 0.54758mV 50147.875p 0.537362mV 50153.623p 0.536322mV 51016.15p 0.548334mV 51086.518p 0.5411mV 51098.9p 0.54018mV 51130.919p 0.535643mV 51169.573p 0.534288mV 52025.571p 0.547911mV 52027.097p 0.547911mV 52035.914p 0.548092mV 52035.947p 0.548092mV 52054.726p 0.549284mV 52072.008p 0.553328mV 52076.693p 0.554709mV 52084.515p 0.55646mV 53056.746p 0.549937mV 53074.921p 0.550136mV 53076.763p 0.550195mV 53082.101p 0.549886mV 53092.128p 0.548161mV 54006.702p 0.54651mV 54007.208p 0.54651mV 54041.473p 0.542858mV 54045.883p 0.542127mV 54066.103p 0.538452mV 55006.134p 0.553519mV 55006.846p 0.553519mV 55018.22p 0.554743mV 55052.056p 0.562548mV 56010.98p 0.552684mV 56011.212p 0.552684mV 56059.753p 0.556589mV 56072.316p 0.557906mV 56109.47p 0.558735mV 57025.309p 0.549961mV 57032.922p 0.548774mV 58005.124p 0.55275mV 58014.288p 0.552327mV 58073.871p 0.556026mV 58088.909p 0.556968mV 58127.203p 0.561023mV 58131.616p 0.56063mV 58142.012p 0.560952mV 59012.27p 0.554942mV 59017.724p 0.555021mV 59023.557p 0.554734mV 59048.648p 0.558789mV 59064.119p 0.561965mV 59064.626p 0.561965mV 59065.03p 0.562784mV 59069.082p 0.562784mV 59087.105p 0.566824mV 60009.458p 0.550707mV 60018.012p 0.550891mV 60021.548p 0.551165mV 61005.406p 0.545687mV 61007.795p 0.545687mV 61018.932p 0.546187mV 61028.725p 0.545221mV 61034.917p 0.54492mV 61054.68p 0.543701mV 61089.12p 0.548076mV 61134.697p 0.557582mV 61134.721p 0.557582mV 61135.05p 0.558355mV 61135.769p 0.558355mV 61139.537p 0.558355mV 61148.348p 0.56027mV 61160.782p 0.561873mV 61161.405p 0.561873mV 61194.724p 0.562562mV 62006.526p 0.548474mV 62008.668p 0.548474mV 62021.977p 0.547008mV 62076.021p 0.540028mV 62110.028p 0.539155mV 62127.779p 0.54014mV 62138.083p 0.540411mV 62141.601p 0.539993mV 63007.462p 0.5502mV 63013.46p 0.549811mV 63051.612p 0.550371mV 63058.117p 0.550352mV 63086.797p 0.549885mV 63093.021p 0.549503mV 63145.274p 0.555611mV 64005.631p 0.550645mV 64027.333p 0.55251mV 64046.425p 0.557308mV 64051.024p 0.55906mV 64063.508p 0.562937mV 65001.567p 0.549359mV 65035.091p 0.552429mV 65038.395p 0.552429mV 66005.105p 0.549551mV 66012.463p 0.549967mV 66054.911p 0.558422mV 66056.16p 0.559211mV 66074.289p 0.559403mV 66078.315p 0.558743mV 66083.126p 0.558452mV 67005.193p 0.55101mV 67050.368p 0.559321mV 68014.773p 0.551491mV 68033.046p 0.555695mV 68033.951p 0.555695mV 69004.027p 0.5477mV 69042.509p 0.548515mV 69055.948p 0.548889mV 69064.092p 0.549254mV 69070.111p 0.551078mV 69114.123p 0.564216mV 69131.595p 0.567913mV 70022.055p 0.549825mV 70025.166p 0.549821mV 70032.462p 0.54945mV 70063.001p 0.544628mV 70071.376p 0.542025mV 71012.146p 0.545117mV 71029.43p 0.546117mV 71040.754p 0.548946mV 71063.207p 0.556145mV 72019.536p 0.554268mV 72059.292p 0.552813mV 72071.613p 0.5509mV 73041.865p 0.555528mV 73052.072p 0.557461mV 73061.957p 0.558667mV 73111.845p 0.556798mV 73117.274p 0.55615mV 73141.409p 0.548194mV 73144.825p 0.548194mV 73181.002p 0.541635mV 73193.341p 0.539992mV 73222.178p 0.532109mV 74037.142p 0.547004mV 74062.946p 0.553976mV 74063.778p 0.553976mV 75005.083p 0.550193mV 75015.425p 0.550642mV 75017.73p 0.550642mV 75036.14p 0.551549mV 75116.235p 0.551697mV 75146.117p 0.549579mV 75147.586p 0.549579mV 75167.04p 0.543333mV 75189.61p 0.534907mV 76059.786p 0.557616mV 76103.529p 0.55804mV 76114.982p 0.556974mV 76158.65p 0.552024mV 76167.044p 0.552425mV 76181.311p 0.553204mV 76184.424p 0.553204mV 76229.708p 0.550414mV 76237.485p 0.548613mV 76250.604p 0.544255mV 76254.987p 0.544255mV 77008.445p 0.548159mV 77012.098p 0.548458mV 77045.216p 0.550536mV 77047.994p 0.550536mV 77081.331p 0.558839mV 77082.982p 0.558839mV 78000.686p 0.551565mV 78002.077p 0.551565mV 78003.446p 0.551565mV 78004.253p 0.551565mV 78045.49p 0.547082mV 78050.163p 0.546045mV 79030.263p 0.552437mV 79048.116p 0.55232mV 79049.717p 0.55232mV 79072.423p 0.551604mV 81008.324p 0.554519mV 81014.613p 0.554187mV 81015.404p 0.554222mV 81020.757p 0.554623mV 81040.962p 0.554775mV 81093.548p 0.553402mV 81127.2p 0.551218mV 81169.935p 0.548771mV 81171.223p 0.54847mV 81179.047p 0.547804mV 81179.708p 0.547804mV 81179.797p 0.547804mV 81184.625p 0.546772mV 81218.137p 0.538094mV 81221.581p 0.53706mV 81257.773p 0.533415mV 81276.588p 0.529912mV 82015.166p 0.548092mV 82033.566p 0.546748mV 82041.474p 0.546458mV 82061.979p 0.546592mV 82064.444p 0.546592mV 82093.144p 0.546379mV 82106.507p 0.546063mV 82168.973p 0.561374mV 83019.675p 0.552622mV 83036.721p 0.556852mV 83057.3p 0.559642mV 83058.599p 0.559642mV 84047.77p 0.553575mV 84061.027p 0.557752mV 85025.107p 0.552157mV 85034.573p 0.551857mV 85036.772p 0.551922mV 85047.165p 0.552419mV 85056.017p 0.553648mV 85074.576p 0.556043mV 85081.617p 0.557279mV 85089.583p 0.557351mV 85125.775p 0.561686mV 87021.67p 0.546662mV 87043.726p 0.542948mV 87054.384p 0.541083mV 87060.738p 0.53848mV 88003.89p 0.549293mV 88018.586p 0.550125mV 88030.271p 0.549872mV 88034.302p 0.549872mV 88062.301p 0.545396mV 88062.715p 0.545396mV 88063.77p 0.545396mV 88114.843p 0.542908mV 88128.5p 0.541643mV 88148.333p 0.534867mV 88148.835p 0.534867mV 89039.417p 0.561003mV 89051.334p 0.566087mV 90008.197p 0.55148mV 90010.745p 0.551871mV 90017.562p 0.551896mV 90039.171p 0.551984mV 90045.014p 0.552388mV 90073.023p 0.551369mV 90103.912p 0.559097mV 90136.088p 0.565394mV 90144.187p 0.567241mV 91004.099p 0.55147mV 91071.306p 0.555486mV 91087.866p 0.550927mV 91088.679p 0.550927mV 91111.95p 0.542108mV 91116.207p 0.540704mV 91122.56p 0.538932mV 93037.343p 0.555877mV 93040.412p 0.556229mV 93042.762p 0.556229mV 93074.99p 0.558032mV 93084.133p 0.557683mV 93089.472p 0.557697mV 93091.628p 0.55808mV 93099.141p 0.558102mV 94017.249p 0.549165mV 94068.996p 0.555553mV 94071.416p 0.555877mV 94078.094p 0.555841mV 94084.133p 0.555444mV 94122.953p 0.549515mV 94154.58p 0.54125mV 94176.112p 0.534179mV 94180.854p 0.533873mV 95005.769p 0.546216mV 95029.079p 0.543937mV 95032.616p 0.542818mV 95033.249p 0.542818mV 95045.5p 0.538724mV 96063.234p 0.548636mV 97001.955p 0.552368mV 97020.529p 0.553265mV 97087.368p 0.557515mV 97111.48p 0.556713mV 97117.944p 0.556045mV 97130.515p 0.555515mV 97161.589p 0.559256mV 97169.429p 0.560801mV 98004.533p 0.547448mV 98005.034p 0.547519mV 98006.979p 0.547519mV 98034.057p 0.544585mV 99011.726p 0.550069mV 99013.984p 0.550069mV 99025.79p 0.546653mV 99027.363p 0.546653mV 99034.201p 0.544783mV 99045.757p 0.537706mV 99054.225p 0.53583mV 100033.939p 0.543722mV 100077.897p 0.536769mV 101070.519p 0.557039mV 101104.737p 0.557665mV 102039.555p 0.552774mV 102048.318p 0.553726mV 102050.877p 0.55475mV 103012.355p 0.550303mV 103013.445p 0.550303mV 103039.766p 0.543494mV 104001.091p 0.551823mV 104036.428p 0.549365mV 104052.296p 0.546913mV 104142.556p 0.546463mV 104147.397p 0.54638mV 104168.349p 0.543858mV 104196.54p 0.539336mV 104196.842p 0.539336mV 104203.846p 0.538883mV 104214.754p 0.53907mV 104231.824p 0.539424mV 104262.721p 0.534786mV 104286.856p 0.532001mV 104287.485p 0.532001mV 104345.015p 0.543206mV 104371.987p 0.550581mV 105001.594p 0.548007mV 105050.052p 0.545514mV 105064.545p 0.544289mV 105093.907p 0.543523mV 106011.154p 0.551774mV 106055.648p 0.555513mV 106059.403p 0.555513mV 106072.551p 0.556777mV 106082.087p 0.558484mV 106090.138p 0.561664mV 107123.193p 0.559098mV 107159.246p 0.552192mV 107195.741p 0.535602mV 108002.836p 0.551583mV 108007.988p 0.551645mV 108053.323p 0.543748mV 108057.142p 0.542331mV 109032.079p 0.554144mV 109037.571p 0.555522mV 110047.736p 0.54938mV 111052.544p 0.552124mV 111059.926p 0.55132mV 112003.295p 0.551874mV 112026.68p 0.552899mV 113001.79p 0.554072mV 113042.117p 0.552816mV 113049.438p 0.553477mV 113056.443p 0.555895mV 114007.528p 0.550712mV 114049.686p 0.553295mV 114080.342p 0.550064mV 114096.229p 0.548444mV 114118.16p 0.54508mV 114118.548p 0.54508mV 114156.623p 0.531759mV 114164.805p 0.529263mV 115023.731p 0.549903mV 115037.703p 0.549267mV 115043.883p 0.54954mV 115045.005p 0.550176mV 115057.942p 0.550346mV 115069.665p 0.549046mV 115088.735p 0.544227mV 116005.018p 0.54967mV 116015.785p 0.550207mV 116023.11p 0.550658mV 116024.226p 0.550658mV 116052.282p 0.547881mV 116056.216p 0.547234mV 116114.022p 0.544336mV 116126.982p 0.545559mV 117007.744p 0.549583mV 117024.034p 0.547605mV 118003.334p 0.549741mV 118007.731p 0.549704mV 118015.602p 0.549997mV 118016.578p 0.549997mV 119022.737p 0.55079mV 119035.291p 0.551339mV 119038.626p 0.551339mV 119045.04p 0.551103mV 119059.076p 0.550874mV 120015.73p 0.549672mV 120026.938p 0.549315mV 120044.782p 0.547122mV 121004.725p 0.552018mV 121005.241p 0.551957mV 121018.096p 0.552935mV 121038.396p 0.557091mV 121054.507p 0.55913mV 121056.127p 0.559815mV 121067.072p 0.561562mV 122008.789p 0.55194mV 122076.355p 0.565308mV 123012.572p 0.553409mV 123020.554p 0.553831mV 123025.41p 0.554593mV 123034.67p 0.554989mV 123048.494p 0.558379mV 124014.799p 0.551642mV 124050.376p 0.542329mV 124052.235p 0.542329mV 124052.461p 0.542329mV 124055.348p 0.542252mV 125012.386p 0.55158mV 125014.345p 0.55158mV 125018.12p 0.552303mV 125024.53p 0.553391mV 125024.992p 0.553391mV 125085.542p 0.561457mV 125093.77p 0.562574mV 126025.95p 0.548624mV 126030.035p 0.548928mV 126062.102p 0.549655mV 126065.948p 0.550326mV 127002.386p 0.55188mV 127033.694p 0.546565mV 127040.503p 0.54454mV 127046.74p 0.542976mV 127047.009p 0.542976mV 127055.723p 0.540934mV 128021.375p 0.545297mV 128022.297p 0.545297mV 128029.552p 0.544578mV 128046.971p 0.538765mV 129029.844p 0.54936mV 129041.152p 0.55177mV 129045.365p 0.553307mV 130011.657p 0.54808mV 130020.437p 0.547553mV 130025.491p 0.54674mV 130032.382p 0.546291mV 130034.958p 0.546291mV 130047.457p 0.547131mV 130078.941p 0.549874mV 130100.872p 0.553427mV 130133.622p 0.55399mV 131010.995p 0.554268mV 131016.706p 0.554193mV 131036.215p 0.551697mV 131037.839p 0.551697mV 131042.724p 0.551254mV 131086.375p 0.556383mV 131105.328p 0.556802mV 131105.752p 0.556802mV 131118.095p 0.558481mV 131135.454p 0.561859mV 132003.485p 0.551727mV 132005.936p 0.551789mV 132016.503p 0.55155mV 132019.41p 0.55155mV 132086.626p 0.557324mV 132120.65p 0.551435mV 132125.225p 0.550812mV 132150.723p 0.547364mV 132162.31p 0.544315mV 132173.2p 0.542003mV 132193.022p 0.536653mV 132218.913p 0.532891mV 132226.783p 0.529116mV 132240.844p 0.522899mV 132242.19p 0.522899mV 133004.181p 0.552329mV 133039.917p 0.545277mV 134041.886p 0.559893mV 134042.79p 0.559893mV 134068.055p 0.563932mV 135063.76p 0.555721mV 135084.61p 0.562674mV 136014.701p 0.548982mV 136027.204p 0.550863mV 136065.782p 0.548896mV 136120.253p 0.528848mV 137016.432p 0.549508mV 137056.737p 0.546688mV 137068.254p 0.544886mV 137077.319p 0.543811mV 138047.757p 0.547295mV 138068.447p 0.549323mV 138082.216p 0.550677mV 138101.286p 0.548369mV 138121.54p 0.543902mV 138160.688p 0.54306mV 138164.777p 0.54306mV 138181.842p 0.543035mV 138184.559p 0.543035mV 138192.644p 0.544864mV 139019.834p 0.550791mV 139047.414p 0.548485mV 139063.923p 0.547895mV 139065.741p 0.547943mV 139116.592p 0.553235mV 139126.338p 0.555198mV 140018.739p 0.547255mV 140060.151p 0.553424mV 140073.576p 0.558013mV 141079.02p 0.546914mV 141107.882p 0.553794mV 141127.509p 0.555201mV 141131.511p 0.555552mV 141132.124p 0.555552mV 141138.981p 0.555538mV 141152.206p 0.555492mV 141166.824p 0.556538mV 141210.519p 0.563268mV 141242.37p 0.578087mV 142004.174p 0.552927mV 142019.504p 0.551808mV 142044.719p 0.549196mV 142050.434p 0.547337mV 143022.979p 0.548476mV 143046.611p 0.544129mV 143047.561p 0.544129mV 143074.315p 0.537185mV 144058.17p 0.548182mV 144092.101p 0.548015mV 144125.724p 0.545926mV 145004.789p 0.550202mV 145027.398p 0.552605mV 146006.816p 0.554377mV 146027.3p 0.553909mV 146064.749p 0.551484mV 146071.312p 0.551997mV 146079.965p 0.55207mV 146107.72p 0.557279mV 146108.499p 0.557279mV 147006.534p 0.552766mV 147008.989p 0.552766mV 147039.896p 0.552609mV 147088.545p 0.54606mV 147094.46p 0.544268mV 147101.218p 0.541046mV 148020.957p 0.547148mV 148045.502p 0.543176mV 148045.922p 0.543176mV 149014.366p 0.553706mV 149022.835p 0.554014mV 149023.74p 0.554014mV 149037.25p 0.555749mV 149041.955p 0.556814mV 149076.503p 0.563555mV 149101.783p 0.567507mV 149104.536p 0.567507mV 150032.578p 0.547043mV 150034.719p 0.547043mV 150035.83p 0.547136mV 150055.002p 0.549709mV 150080.125p 0.554237mV 150095.689p 0.555672mV 150099.675p 0.555672mV 150113.418p 0.556779mV 150113.984p 0.556779mV 150114.326p 0.556779mV 151033.17p 0.557565mV 151036.18p 0.557519mV 151045.22p 0.55853mV 151047.655p 0.55853mV 152000.506p 0.553992mV 152011.571p 0.553783mV 152020.315p 0.554301mV 152021.147p 0.554301mV 153036.087p 0.560228mV 154026.19p 0.546802mV 154036.7p 0.547164mV 154040.228p 0.547527mV 154062.698p 0.547502mV 154063.86p 0.547502mV 154097.649p 0.547039mV 154110.942p 0.544774mV 155036.578p 0.550162mV 155041.296p 0.549844mV 156065.513p 0.554523mV 156083.777p 0.558134mV 157036.311p 0.542454mV 158002.291p 0.552143mV 158012.039p 0.551727mV 158034.481p 0.547219mV 158040.649p 0.544585mV 158042.753p 0.544585mV 158048.939p 0.543081mV 158049.569p 0.543081mV 159027.958p 0.551386mV 159036.141p 0.552503mV 159047.233p 0.555093mV 160021.088p 0.552165mV 160026.678p 0.551427mV 160039.11p 0.550317mV 160078.0p 0.547281mV 160106.77p 0.54307mV 161038.87p 0.549918mV 161058.957p 0.548871mV 161063.915p 0.548426mV 161064.52p 0.548426mV 161086.407p 0.548022mV 161164.479p 0.556974mV 161178.54p 0.555656mV 161183.935p 0.555223mV 161186.293p 0.554427mV 161193.133p 0.553269mV 161204.615p 0.550592mV 161238.386p 0.535212mV 162034.661p 0.546384mV 162043.544p 0.547659mV 162055.954p 0.549026mV 162059.793p 0.549026mV 162072.362p 0.551495mV 163000.044p 0.547713mV 163005.31p 0.547643mV 163007.008p 0.547643mV 164004.402p 0.551771mV 164024.386p 0.554107mV 164032.457p 0.555284mV 164053.008p 0.558397mV 165017.749p 0.546787mV 165041.082p 0.551022mV 167046.556p 0.53669mV 168001.799p 0.549174mV 168004.845p 0.549174mV 168006.37p 0.54919mV 168007.266p 0.54919mV 168047.976p 0.555195mV 168051.251p 0.555588mV 168053.404p 0.555588mV 168065.996p 0.557516mV 169007.265p 0.547069mV 169058.567p 0.553037mV 169061.2p 0.553382mV 169084.786p 0.553316mV 169086.498p 0.554035mV 169103.778p 0.556207mV 169137.684p 0.555915mV 169144.258p 0.556307mV 170003.046p 0.553533mV 170020.423p 0.553155mV 170059.091p 0.558684mV 171049.939p 0.561168mV 172005.141p 0.548529mV 172016.977p 0.548001mV 172024.065p 0.548287mV 172038.758p 0.548417mV 172054.494p 0.549653mV 172071.583p 0.54937mV 172095.597p 0.553451mV 173011.002p 0.547974mV 173014.978p 0.547974mV 173024.487p 0.54767mV 173033.314p 0.546635mV 173054.683p 0.54896mV 173070.604p 0.554222mV 173076.958p 0.556456mV 174025.577p 0.547708mV 174027.097p 0.547708mV 174078.98p 0.549807mV 174102.136p 0.552185mV 174108.818p 0.553033mV 174109.204p 0.553033mV 174129.246p 0.552811mV 174154.813p 0.548063mV 174159.613p 0.54676mV 174178.727p 0.543778mV 174191.097p 0.542129mV 174202.146p 0.540686mV 174204.154p 0.540686mV 175045.011p 0.557966mV 175048.159p 0.557966mV 176046.851p 0.542459mV 176051.668p 0.541405mV 177032.42p 0.551061mV 178000.336p 0.546306mV 178031.054p 0.546366mV 178050.21p 0.551795mV 178052.255p 0.551795mV 179001.361p 0.549073mV 179038.593p 0.542432mV 179047.869p 0.538278mV 180018.728p 0.552532mV 180060.217p 0.551441mV 180076.139p 0.550566mV 180119.85p 0.549576mV 181008.485p 0.547759mV 181028.533p 0.548548mV 181043.474p 0.550782mV 181065.015p 0.553784mV 181078.261p 0.554192mV 181136.555p 0.542138mV 182025.767p 0.550851mV 182033.434p 0.549831mV 182044.95p 0.547419mV 182053.525p 0.545727mV 183007.592p 0.546442mV 183038.45p 0.548242mV 183053.859p 0.547494mV 183072.258p 0.546737mV 183073.792p 0.546737mV 183085.09p 0.544149mV 183101.671p 0.543375mV 183106.92p 0.543356mV 183108.101p 0.543356mV 183114.921p 0.5437mV 183174.572p 0.562306mV 183179.165p 0.564468mV 184005.314p 0.550962mV 184043.203p 0.550111mV 184048.123p 0.549367mV 184154.195p 0.55087mV 184159.312p 0.552315mV 185001.808p 0.552594mV 185017.772p 0.553432mV 186007.125p 0.552504mV 186009.947p 0.552504mV 186024.205p 0.552729mV 187001.764p 0.546042mV 187002.645p 0.546042mV 187017.296p 0.545191mV 187023.749p 0.544909mV 187059.885p 0.537809mV 188014.75p 0.552548mV 189001.172p 0.547783mV 189047.261p 0.552517mV 189053.419p 0.55366mV 189054.844p 0.55366mV 189055.186p 0.555173mV 190128.209p 0.556125mV 191017.292p 0.547322mV 191028.332p 0.549783mV 192012.253p 0.5499mV 192012.874p 0.5499mV 192025.681p 0.550356mV 192043.181p 0.550461mV 192051.313p 0.551636mV 192057.752p 0.551678mV 192088.739p 0.550889mV 192096.52p 0.55065mV 192115.824p 0.550211mV 192117.61p 0.550211mV 193013.566p 0.547946mV 194009.317p 0.552542mV 194019.903p 0.551565mV 195006.179p 0.549615mV 195029.747p 0.545843mV 195032.059p 0.544718mV 195033.85p 0.544718mV 195039.609p 0.543959mV 195042.595p 0.543566mV 195048.377p 0.542805mV 195100.232p 0.535765mV 196011.287p 0.550606mV 196034.301p 0.553901mV 196046.93p 0.556753mV 196047.627p 0.556753mV 196070.747p 0.560589mV 196070.782p 0.560589mV 197001.045p 0.547645mV 197004.897p 0.547645mV 197008.826p 0.547676mV 197022.384p 0.549238mV 197032.328p 0.548943mV 197036.401p 0.548981mV 197057.019p 0.552074mV 197066.832p 0.552536mV 197072.662p 0.552224mV 197076.861p 0.551549mV 197077.963p 0.551549mV 197110.811p 0.550572mV 198004.613p 0.549132mV 198052.631p 0.542977mV 198079.42p 0.542608mV 198111.224p 0.537625mV 199006.182p 0.552913mV 199019.632p 0.553993mV 199067.909p 0.553602mV 200003.656p 0.55087mV 200004.061p 0.55087mV 200089.819p 0.559155mV 201006.92p 0.552516mV 201007.091p 0.552516mV 201010.103p 0.552831mV 201015.704p 0.552778mV 201021.489p 0.552359mV 201037.776p 0.548899mV 202010.735p 0.553619mV 202031.221p 0.553595mV 202036.149p 0.554321mV 202039.096p 0.554321mV 202042.854p 0.555413mV 202043.551p 0.555413mV 202044.305p 0.555413mV 202082.843p 0.563478mV 203002.077p 0.553877mV 203006.112p 0.553834mV 203027.987p 0.553648mV 203063.158p 0.549602mV 204001.966p 0.546469mV 204042.665p 0.553203mV 205000.48p 0.553287mV 205025.88p 0.551429mV 205041.383p 0.549738mV 206020.26p 0.550558mV 206059.834p 0.552513mV 206080.838p 0.555383mV 206119.76p 0.560371mV 207003.216p 0.546952mV 207008.653p 0.547015mV 207033.906p 0.546216mV 207038.522p 0.545541mV 207055.224p 0.545018mV 207066.723p 0.544012mV 207068.292p 0.544012mV 207071.053p 0.543688mV 208001.837p 0.552938mV 208070.483p 0.54855mV 208077.117p 0.547173mV 208095.148p 0.54239mV 208097.046p 0.54239mV 208099.556p 0.54239mV 209012.435p 0.551365mV 209012.873p 0.551365mV 209036.511p 0.550884mV 209039.494p 0.550884mV 209054.14p 0.551755mV 209056.157p 0.552531mV 209056.88p 0.552531mV 209067.397p 0.552983mV 209083.915p 0.555304mV 210017.406p 0.550444mV 210022.713p 0.550785mV 210024.062p 0.550785mV 210026.059p 0.551491mV 210043.305p 0.552141mV 210124.232p 0.557549mV 210149.361p 0.560365mV 210150.309p 0.560713mV 210165.327p 0.5625mV 210191.085p 0.562118mV 210198.135p 0.562124mV 210198.447p 0.562124mV 210214.407p 0.562159mV 210222.889p 0.564025mV 211019.695p 0.552995mV 211019.959p 0.552995mV 211077.582p 0.553042mV 211084.154p 0.552627mV 211095.333p 0.551393mV 211118.48p 0.549769mV 211119.555p 0.549769mV 211138.899p 0.551096mV 212003.574p 0.554459mV 212035.956p 0.549602mV 212045.02p 0.549401mV 213002.654p 0.548432mV 213023.646p 0.549054mV 213032.886p 0.550104mV 214025.479p 0.551472mV 215003.997p 0.553555mV 215029.958p 0.554987mV 215075.626p 0.559735mV 215078.97p 0.559735mV 215084.0p 0.560111mV 215088.959p 0.560124mV 215099.751p 0.560525mV 215105.538p 0.560207mV 215111.431p 0.559872mV 215162.098p 0.554895mV 216005.53p 0.550444mV 216007.189p 0.550444mV 216020.71p 0.549494mV 216031.819p 0.548256mV 216093.675p 0.53863mV 216108.636p 0.535828mV 216115.375p 0.533092mV 217003.88p 0.5527mV 217089.473p 0.560664mV 217111.64p 0.563728mV 217113.069p 0.563728mV 218033.153p 0.548501mV 218064.846p 0.540023mV 218079.068p 0.535209mV 219008.224p 0.550728mV 219019.993p 0.551275mV 219033.111p 0.553734mV 219077.677p 0.565536mV 219080.906p 0.566739mV 220001.946p 0.546397mV 220016.209p 0.546941mV 220019.913p 0.546941mV 220050.342p 0.548855mV 220056.615p 0.548926mV 220065.691p 0.549438mV 220066.578p 0.549438mV 220075.12p 0.548497mV 220102.939p 0.543441mV 220107.642p 0.541338mV 220126.569p 0.533658mV 220135.572p 0.52981mV 220140.575p 0.527334mV 221010.532p 0.55314mV 221011.49p 0.55314mV 221012.099p 0.55314mV 221013.591p 0.55314mV 221020.094p 0.552895mV 221070.708p 0.556783mV 221071.74p 0.556783mV 221091.963p 0.554843mV 221120.939p 0.557067mV 221121.837p 0.557067mV 221124.39p 0.557067mV 221135.834p 0.556176mV 221138.211p 0.556176mV 221141.683p 0.555881mV 221146.844p 0.555221mV 221150.822p 0.554927mV 221208.947p 0.555374mV 221209.609p 0.555374mV 223006.965p 0.548356mV 223017.358p 0.547175mV 223024.244p 0.546037mV 223039.015p 0.542628mV 223063.529p 0.54059mV 224003.247p 0.551461mV 224007.211p 0.551481mV 224024.859p 0.552281mV 225011.512p 0.554729mV 225056.187p 0.559369mV 226034.283p 0.545325mV 226055.212p 0.540962mV 227017.521p 0.553508mV 227027.773p 0.55442mV 227028.511p 0.55442mV 227055.549p 0.557145mV 227068.02p 0.557323mV 227086.274p 0.557684mV 227101.308p 0.560339mV 227107.286p 0.561714mV 227115.032p 0.564836mV 228005.566p 0.550072mV 228050.947p 0.553525mV 228079.28p 0.557666mV 229024.152p 0.549387mV 229061.417p 0.550501mV 229071.557p 0.550244mV 229085.044p 0.547126mV 229099.624p 0.545418mV 230013.506p 0.546735mV 230034.008p 0.54864mV 230051.198p 0.549812mV 230052.779p 0.549812mV 230067.76p 0.549234mV 230079.587p 0.54873mV 230092.403p 0.546332mV 230112.657p 0.543133mV 230118.235p 0.543062mV 230132.148p 0.545034mV 230144.795p 0.548172mV 230145.088p 0.549558mV 230157.268p 0.551966mV 230173.869p 0.553944mV 230188.658p 0.55485mV 230203.045p 0.554691mV 231011.722p 0.551856mV 231032.962p 0.549705mV 231043.48p 0.54789mV 231050.06p 0.546068mV 232008.794p 0.547854mV 232038.181p 0.553851mV 232046.656p 0.557083mV 233002.62p 0.550001mV 233029.274p 0.550354mV 233035.38p 0.551595mV 233042.849p 0.552033mV 233044.692p 0.552033mV 233064.455p 0.557457mV 234011.944p 0.55277mV 234023.626p 0.553247mV 234026.488p 0.553301mV 234078.465p 0.557094mV 234078.942p 0.557094mV 234083.952p 0.556776mV 234087.87p 0.556824mV 234108.153p 0.559942mV 234129.433p 0.5638mV 234135.966p 0.5672mV 235019.252p 0.54793mV 235028.013p 0.549073mV 235028.579p 0.549073mV 235034.406p 0.549462mV 235046.195p 0.548441mV 235057.318p 0.545937mV 236010.204p 0.552604mV 236021.932p 0.552128mV 236028.726p 0.55134mV 236044.93p 0.550436mV 236065.033p 0.55086mV 237009.995p 0.552999mV 237012.468p 0.552637mV 237027.217p 0.552273mV 237028.021p 0.552273mV 237038.585p 0.55117mV 237054.633p 0.549683mV 237069.31p 0.550732mV 237076.55p 0.55178mV 237088.215p 0.554279mV 237093.295p 0.555341mV 237114.493p 0.558106mV 237137.344p 0.560053mV 237158.391p 0.559078mV 238006.492p 0.551407mV 238008.048p 0.551407mV 238053.479p 0.551326mV 238086.279p 0.557113mV 239026.863p 0.54483mV 239047.063p 0.540338mV 239053.601p 0.53848mV 239061.423p 0.534392mV 240008.967p 0.553516mV 240024.238p 0.553582mV 240043.985p 0.557329mV 240094.069p 0.55876mV 240095.951p 0.558806mV 240098.094p 0.558806mV 240111.676p 0.557501mV 240118.988p 0.557559mV 240146.467p 0.558345mV 240148.411p 0.558345mV 241029.772p 0.553882mV 241069.403p 0.555521mV 241091.959p 0.557015mV 241096.812p 0.556952mV 241120.113p 0.562154mV 242012.425p 0.553668mV 242029.243p 0.556058mV 242058.61p 0.558298mV 242098.678p 0.560178mV 242105.96p 0.560498mV 242108.352p 0.560498mV 242114.568p 0.560116mV 242150.132p 0.552845mV 242151.774p 0.552845mV 243005.082p 0.552405mV 243013.902p 0.552728mV 243035.63p 0.553989mV 243050.255p 0.55681mV 243054.25p 0.55681mV 244017.159p 0.54729mV 244038.507p 0.553302mV 244065.324p 0.556874mV 244066.464p 0.556874mV 244094.252p 0.553903mV 244109.075p 0.553032mV 244112.367p 0.553478mV 245017.981p 0.551915mV 245020.179p 0.550836mV 245077.296p 0.54617mV 245087.646p 0.545054mV 245091.74p 0.544673mV 246001.059p 0.553307mV 246007.04p 0.553343mV 246035.779p 0.550249mV 246047.294p 0.548475mV 246050.811p 0.548133mV 246061.609p 0.546342mV 247007.069p 0.549442mV 247011.999p 0.549784mV 247019.818p 0.54976mV 247043.862p 0.548523mV 247069.718p 0.546879mV 247074.257p 0.54647mV 248002.625p 0.554674mV 248012.339p 0.555128mV 249000.362p 0.549817mV 249009.756p 0.54974mV 249013.845p 0.549297mV 249022.044p 0.548043mV 249037.631p 0.544507mV 249047.361p 0.541043mV 250009.379p 0.553447mV 250017.497p 0.553817mV 250057.739p 0.555991mV 250115.796p 0.562558mV 250123.902p 0.562933mV 250136.325p 0.564074mV 250141.718p 0.563731mV 250158.333p 0.562721mV 250172.2p 0.56211mV 250190.849p 0.559402mV 250244.394p 0.547444mV 251011.433p 0.546268mV 251024.54p 0.546652mV 251027.802p 0.547396mV 251045.79p 0.54673mV 251105.08p 0.5383mV 251126.718p 0.533309mV 251139.751p 0.529346mV 251148.81p 0.523913mV 252016.315p 0.545822mV 252044.472p 0.544357mV 252056.446p 0.544209mV 253018.989p 0.550849mV 253021.134p 0.549695mV 253050.187p 0.549706mV 253050.245p 0.549706mV 253060.037p 0.549947mV 253074.395p 0.55165mV 253079.819p 0.55305mV 253097.123p 0.559391mV 253101.251p 0.560433mV 254003.834p 0.553006mV 254007.059p 0.552916mV 254032.077p 0.552102mV 254041.673p 0.551556mV 254102.765p 0.54461mV 254115.198p 0.54029mV 254120.798p 0.539088mV 255019.88p 0.553329mV 255020.326p 0.552937mV 255032.446p 0.551784mV 255035.107p 0.551023mV 255041.64p 0.550626mV 255060.792p 0.548289mV 255077.333p 0.546325mV 255086.297p 0.545119mV 256014.798p 0.554121mV 256020.168p 0.553659mV 256049.173p 0.552677mV 256087.975p 0.5522mV 256123.065p 0.552396mV 256186.78p 0.576624mV 256186.857p 0.576624mV 256192.097p 0.580533mV 256199.595p 0.584809mV 257069.98p 0.565084mV 258000.121p 0.546705mV 258023.815p 0.545386mV 258072.162p 0.540118mV 259007.725p 0.546344mV 259046.811p 0.544459mV 259047.224p 0.544459mV 259068.331p 0.542802mV 259068.648p 0.542802mV 259071.811p 0.542389mV 259136.146p 0.539598mV 259154.303p 0.540195mV 259184.881p 0.543247mV 260039.545p 0.562521mV 261030.001p 0.551558mV 261036.684p 0.551611mV 261044.326p 0.551297mV 261064.626p 0.55003mV 261071.528p 0.549753mV 261081.535p 0.548006mV 261083.213p 0.548006mV 262001.023p 0.545938mV 262007.537p 0.545967mV 262007.602p 0.545967mV 262011.269p 0.546362mV 262014.579p 0.546362mV 262034.7p 0.549403mV 262086.882p 0.542841mV 262099.228p 0.540353mV 262108.542p 0.537127mV 262115.531p 0.533159mV 263016.537p 0.554721mV 263020.554p 0.55501mV 263022.23p 0.55501mV 263025.884p 0.554933mV 263036.633p 0.554416mV 263072.977p 0.553892mV 263086.774p 0.553305mV 263094.583p 0.553597mV 263131.51p 0.563275mV 264045.538p 0.547046mV 264053.746p 0.547378mV 264073.659p 0.549415mV 264116.755p 0.558471mV 264148.642p 0.562917mV 264177.963p 0.566657mV 264179.203p 0.566657mV 264200.504p 0.569739mV 264208.0p 0.570433mV 264217.048p 0.572924mV 264217.643p 0.572924mV 264217.856p 0.572924mV 265023.994p 0.551867mV 265070.768p 0.541326mV 265073.36p 0.541326mV 265090.481p 0.539095mV 266004.014p 0.552613mV 266011.977p 0.552913mV 266030.104p 0.557188mV 266053.575p 0.559312mV 267022.39p 0.548423mV 267066.842p 0.539261mV 268016.611p 0.550701mV 268019.769p 0.550701mV 268027.314p 0.550148mV 268034.276p 0.549687mV 268084.508p 0.55196mV 268085.904p 0.551852mV 268107.654p 0.549949mV 268161.674p 0.55663mV 268170.824p 0.557457mV 268179.245p 0.558052mV 268188.027p 0.558141mV 268210.648p 0.557058mV 268214.536p 0.557058mV 269073.439p 0.546755mV 269089.833p 0.550196mV 269099.996p 0.552861mV 269103.169p 0.554014mV 270005.965p 0.553183mV 271029.157p 0.547681mV 271029.486p 0.547681mV 271054.676p 0.544343mV 272011.112p 0.55221mV 272057.687p 0.552486mV 272074.007p 0.55454mV 272077.655p 0.555958mV 272095.052p 0.559459mV 272101.233p 0.559794mV 272113.852p 0.559382mV 272134.735p 0.557882mV 272139.063p 0.557154mV 272143.536p 0.556796mV 273005.845p 0.54781mV 273051.851p 0.550388mV 273062.222p 0.552058mV 273067.781p 0.553442mV 273087.731p 0.556797mV 274006.084p 0.549472mV 274037.386p 0.543128mV 274044.332p 0.541277mV 275024.7p 0.549294mV 275106.273p 0.545558mV 276004.845p 0.545949mV 276007.066p 0.546029mV 276014.101p 0.546474mV 276018.551p 0.547283mV 276018.615p 0.547283mV 276027.102p 0.5478mV 276057.954p 0.544212mV 276062.216p 0.543183mV 276067.906p 0.541785mV 276072.11p 0.540019mV 277079.158p 0.555879mV 278013.36p 0.553331mV 278034.913p 0.548583mV 278055.943p 0.543705mV 279001.711p 0.551512mV 279060.925p 0.558553mV 279063.996p 0.558553mV 280078.334p 0.550874mV 280087.712p 0.548227mV 281013.626p 0.546616mV 281018.347p 0.54741mV 281069.053p 0.550607mV 281081.191p 0.551548mV 281112.17p 0.55531mV 281126.665p 0.554492mV 281132.669p 0.553496mV 281135.561p 0.55287mV 281165.53p 0.546625mV 281177.273p 0.545056mV 281209.997p 0.543344mV 282000.329p 0.552648mV 282017.975p 0.553808mV 282047.751p 0.555802mV 282061.176p 0.558109mV 282065.812p 0.559615mV 282067.287p 0.559615mV 282071.323p 0.561489mV 283011.688p 0.545135mV 283018.666p 0.545094mV 283026.902p 0.543914mV 283032.565p 0.543506mV 283048.58p 0.541545mV 283050.587p 0.540401mV 283053.86p 0.540401mV 283060.978p 0.537742mV 283065.967p 0.536225mV 283070.257p 0.534341mV 284049.142p 0.541726mV 284054.228p 0.540627mV 284068.187p 0.536592mV 285008.1p 0.547918mV 285022.562p 0.548548mV 285022.611p 0.548548mV 285027.009p 0.548512mV 285033.601p 0.548109mV 285046.897p 0.546894mV 285094.968p 0.542405mV 285098.41p 0.540876mV 286000.92p 0.549105mV 286025.378p 0.550978mV 286086.334p 0.559209mV 287017.648p 0.547705mV 287037.527p 0.549977mV 287068.868p 0.552687mV 287079.199p 0.553847mV 288031.97p 0.552369mV 288048.844p 0.551274mV 288067.051p 0.546903mV 288070.61p 0.545811mV 288075.414p 0.544352mV 288088.189p 0.541066mV 288092.482p 0.539238mV 288096.921p 0.537773mV 288105.3p 0.535199mV 289011.224p 0.546673mV 289037.744p 0.547994mV 289057.462p 0.547893mV 289095.188p 0.543349mV 289152.466p 0.542436mV 289172.437p 0.543114mV 289181.172p 0.542729mV 289222.434p 0.54419mV 290001.387p 0.547642mV 290003.713p 0.547642mV 290007.448p 0.547621mV 290032.716p 0.548617mV 290034.386p 0.548617mV 290046.502p 0.551857mV 290057.679p 0.55439mV 290067.787p 0.556204mV 290070.068p 0.556568mV 291012.782p 0.553045mV 291016.369p 0.553806mV 291040.007p 0.558699mV 291057.794p 0.562081mV 291067.909p 0.563249mV 292005.336p 0.547538mV 292009.581p 0.547538mV 292025.48p 0.549979mV 292051.194p 0.555793mV 292051.541p 0.555793mV 292052.885p 0.555793mV 293023.86p 0.543339mV 293039.74p 0.539414mV 293047.704p 0.535449mV 293058.836p 0.532206mV 294007.954p 0.548486mV 295031.375p 0.551258mV 296024.699p 0.55041mV 296028.505p 0.551141mV 296051.853p 0.552993mV 296052.09p 0.552993mV 296068.294p 0.554133mV 297034.2p 0.542514mV 297041.182p 0.539824mV 298042.293p 0.552554mV 298080.174p 0.555959mV 298108.367p 0.559208mV 298163.988p 0.560868mV 298167.643p 0.560243mV 298191.417p 0.558273mV 298201.578p 0.555982mV 298238.577p 0.544261mV 298245.913p 0.539117mV 299023.222p 0.552202mV 299054.747p 0.552822mV 299060.777p 0.554742mV 299071.466p 0.556667mV 300007.415p 0.550772mV 300028.835p 0.549291mV 300040.056p 0.546348mV 300047.293p 0.545609mV 300069.171p 0.542631mV 300090.902p 0.542125mV 300091.101p 0.542125mV 301003.949p 0.550208mV 301065.288p 0.542532mV 302013.076p 0.545488mV 302037.192p 0.541498mV 302038.365p 0.541498mV 303010.497p 0.552638mV 303043.19p 0.550501mV 303049.485p 0.551303mV 303076.678p 0.554284mV 303078.254p 0.554284mV 303092.24p 0.554502mV 303096.011p 0.554577mV 303096.668p 0.554577mV 303118.248p 0.556353mV 303119.852p 0.556353mV 303130.506p 0.558799mV 304048.362p 0.537421mV 305031.721p 0.556756mV 305037.625p 0.5574mV 306010.36p 0.55142mV 306036.34p 0.551465mV 306062.661p 0.546048mV 306089.92p 0.54245mV 306111.197p 0.540634mV 306114.097p 0.540634mV 306150.06p 0.554421mV 307014.785p 0.548601mV 307038.343p 0.549288mV 307070.316p 0.54854mV 307070.454p 0.54854mV 307092.434p 0.551484mV 308006.373p 0.54708mV 308011.605p 0.547395mV 308017.438p 0.548077mV 308034.042p 0.550124mV 309004.472p 0.547095mV 309023.087p 0.547136mV 309029.009p 0.547881mV 309051.816p 0.54833mV 309083.742p 0.545926mV 309096.294p 0.545656mV 309125.699p 0.54041mV 309131.977p 0.539358mV 309143.71p 0.536158mV 309174.698p 0.528748mV 309178.568p 0.527325mV 309178.623p 0.527325mV 310011.958p 0.547007mV 310015.89p 0.547036mV 310063.911p 0.555718mV 310077.159p 0.557667mV 312022.772p 0.550092mV 312024.102p 0.550092mV 312032.079p 0.548254mV 312037.766p 0.547516mV 312059.57p 0.545271mV 312096.675p 0.550851mV 312112.47p 0.557277mV 312128.776p 0.564788mV 312141.707p 0.572668mV 312147.212p 0.575543mV 313035.046p 0.549665mV 313067.974p 0.553142mV 313075.947p 0.552849mV 313094.802p 0.552969mV 313112.925p 0.550224mV 313116.298p 0.54881mV 313119.808p 0.54881mV 313130.98p 0.545299mV 313182.899p 0.543885mV 313221.61p 0.537512mV 314010.167p 0.546439mV 314014.278p 0.546439mV 314022.661p 0.545179mV 314060.707p 0.538605mV 315033.595p 0.558147mV 315034.211p 0.558147mV 315042.089p 0.559297mV 315049.226p 0.559329mV 315050.899p 0.558999mV 315052.767p 0.558999mV 315053.494p 0.558999mV 315054.387p 0.558999mV 315098.662p 0.549983mV 316012.843p 0.54763mV 316037.268p 0.550362mV 316052.211p 0.550239mV 316055.348p 0.550199mV 317004.959p 0.550505mV 317005.771p 0.550435mV 317020.722p 0.548762mV 317042.215p 0.548481mV 317073.593p 0.538902mV 318002.656p 0.552641mV 318010.999p 0.552118mV 319007.401p 0.552289mV 319009.439p 0.552289mV 319009.879p 0.552289mV 319025.124p 0.550971mV 319032.564p 0.551371mV 319039.978p 0.551403mV 319043.549p 0.551068mV 319055.674p 0.552249mV 319088.728p 0.56007mV 320012.75p 0.545721mV 320016.095p 0.545707mV 320023.416p 0.546059mV 320025.808p 0.546776mV 320059.257p 0.554377mV 321010.325p 0.552121mV 321059.891p 0.546096mV 321076.582p 0.539425mV 322018.17p 0.553231mV 322026.155p 0.552036mV 322047.264p 0.545969mV 322047.684p 0.545969mV 323038.182p 0.549428mV 323043.763p 0.548303mV 324019.017p 0.54567mV 324039.19p 0.547342mV 324067.933p 0.545088mV 324093.758p 0.543484mV 324100.64p 0.543922mV 324131.542p 0.543704mV 325032.633p 0.545009mV 325038.604p 0.544937mV 325042.774p 0.545229mV 325051.573p 0.545443mV 325051.879p 0.545443mV 325080.083p 0.547511mV 325113.94p 0.547336mV 325117.294p 0.54724mV 325119.733p 0.54724mV 325126.83p 0.546675mV 325141.791p 0.54855mV 325157.383p 0.552959mV 325167.607p 0.556009mV 325208.387p 0.558658mV 326014.011p 0.553904mV 326014.295p 0.553904mV 326025.507p 0.55379mV 326053.435p 0.553835mV 326081.28p 0.549541mV 327031.493p 0.542016mV 327034.076p 0.542016mV 327046.139p 0.540216mV 327087.02p 0.546099mV 327089.949p 0.546099mV 328005.72p 0.548041mV 328008.397p 0.548041mV 328031.108p 0.54787mV 328042.388p 0.549771mV 328059.182p 0.551705mV 328091.163p 0.55782mV 328091.412p 0.55782mV 328099.757p 0.559326mV 328101.504p 0.560469mV 328101.8p 0.560469mV 328112.041p 0.56386mV 329001.419p 0.545477mV 329002.563p 0.545477mV 329018.716p 0.546845mV 329020.267p 0.547302mV 329040.081p 0.546948mV 329095.044p 0.546285mV 329106.613p 0.543964mV 329109.731p 0.543964mV 329137.428p 0.537761mV 329158.563p 0.530215mV 329164.884p 0.527777mV 329165.016p 0.524971mV 330004.945p 0.55136mV 330005.814p 0.551432mV 330039.45p 0.547832mV 330046.998p 0.546867mV 330087.025p 0.545094mV 330180.131p 0.578033mV 330186.477p 0.580936mV 330202.135p 0.588925mV 330209.769p 0.591838mV 331009.403p 0.547633mV 331032.27p 0.544669mV 331035.716p 0.543857mV 331058.318p 0.538407mV 331062.277p 0.536491mV 332022.543p 0.55022mV 332024.419p 0.55022mV 332041.97p 0.547028mV 332087.973p 0.544234mV 332089.958p 0.544234mV 332097.279p 0.54446mV 332113.128p 0.544246mV 332153.035p 0.536326mV 333000.327p 0.546366mV 333022.473p 0.548869mV 333054.642p 0.557769mV 334045.795p 0.549219mV 334051.097p 0.549623mV 334068.842p 0.551563mV 334074.793p 0.552697mV 334079.132p 0.553466mV 334080.416p 0.55387mV 334086.828p 0.55464mV 334087.059p 0.55464mV 334115.797p 0.563313mV 334119.692p 0.563313mV 335046.969p 0.545741mV 336032.677p 0.547236mV 336037.944p 0.545793mV 336051.47p 0.54072mV 337044.77p 0.54867mV 337070.044p 0.544109mV 337082.365p 0.543076mV 337090.647p 0.542771mV 337104.414p 0.543192mV 337116.718p 0.545094mV 337133.376p 0.545161mV 337136.224p 0.545183mV 337156.073p 0.542339mV 337164.713p 0.541991mV 337185.655p 0.542053mV 337206.227p 0.539138mV 338044.677p 0.547392mV 338090.578p 0.546338mV 338124.027p 0.547838mV 338136.389p 0.545458mV 339005.43p 0.545672mV 339059.733p 0.550526mV 339069.372p 0.551669mV 340017.361p 0.546225mV 340048.85p 0.542128mV 341006.276p 0.549979mV 341006.854p 0.549979mV 341082.859p 0.56314mV 342034.851p 0.550425mV 343016.556p 0.550338mV 343024.758p 0.54991mV 343066.918p 0.54636mV 343092.171p 0.549228mV 343121.636p 0.547565mV 344020.845p 0.548619mV 344036.945p 0.548013mV 344077.963p 0.550263mV 344084.767p 0.551271mV 344093.497p 0.553655mV 345003.96p 0.55071mV 345028.572p 0.550254mV 345051.184p 0.541409mV 346027.399p 0.550101mV 346030.032p 0.551201mV 346033.028p 0.551201mV 346041.169p 0.553764mV 346049.62p 0.554497mV 347075.234p 0.553309mV 347084.82p 0.55366mV 347119.244p 0.56129mV 348005.54p 0.551377mV 348006.948p 0.551377mV 348034.115p 0.553635mV 348057.623p 0.558453mV 348061.615p 0.559638mV 348105.782p 0.562001mV 348113.094p 0.562481mV 349003.113p 0.545425mV 349022.457p 0.547262mV 349052.158p 0.555911mV 350005.897p 0.552824mV 350006.08p 0.552824mV 350007.268p 0.552824mV 350008.124p 0.552824mV 350045.417p 0.552875mV 350045.702p 0.552875mV 350066.906p 0.555477mV 350067.219p 0.555477mV 350099.917p 0.559803mV 350100.743p 0.560109mV 350107.688p 0.560055mV 351030.091p 0.555319mV 352015.052p 0.552296mV 352032.739p 0.552386mV 352035.719p 0.552419mV 352043.483p 0.552818mV 352063.03p 0.553695mV 352068.682p 0.554467mV 352074.803p 0.554875mV 352088.196p 0.556113mV 352090.319p 0.5558mV 352106.992p 0.552691mV 352109.665p 0.552691mV 352128.78p 0.548586mV 352130.055p 0.546834mV 352134.639p 0.546834mV 352137.833p 0.544719mV 352146.674p 0.540857mV 352150.386p 0.538379mV 352175.132p 0.527071mV 353020.242p 0.549786mV 353028.273p 0.550519mV 353034.153p 0.550888mV 353036.675p 0.550894mV 353053.797p 0.551659mV 353055.663p 0.551677mV 353065.83p 0.552088mV 353088.62p 0.548573mV 353126.825p 0.542456mV 353141.809p 0.539767mV 353156.25p 0.536022mV 354002.041p 0.54862mV 354018.428p 0.549225mV 354021.658p 0.549674mV 354021.857p 0.549674mV 354046.564p 0.550107mV 354068.196p 0.546825mV 354123.7p 0.534719mV 355014.502p 0.553901mV 355023.866p 0.552853mV 355053.292p 0.556253mV 355137.857p 0.557718mV 355142.425p 0.558791mV 355143.635p 0.558791mV 355171.148p 0.557494mV 356049.353p 0.552495mV 357005.118p 0.548497mV 357050.105p 0.543271mV 357073.854p 0.538258mV 357074.782p 0.538258mV 358009.911p 0.552605mV 358033.712p 0.549696mV 358036.23p 0.54831mV 358051.35p 0.541951mV 359017.708p 0.546194mV 359045.787p 0.544534mV 359045.824p 0.544534mV 360047.467p 0.559311mV 361040.779p 0.540273mV 361044.761p 0.540273mV 362013.561p 0.552057mV 362019.4p 0.551988mV 362033.744p 0.549578mV 362037.339p 0.548041mV 363009.064p 0.548338mV 363052.077p 0.550336mV 363075.334p 0.550754mV 363081.912p 0.551059mV 363082.031p 0.551059mV 363103.769p 0.550094mV 363122.108p 0.547676mV 363151.719p 0.541848mV 363163.898p 0.542087mV 363172.301p 0.54378mV 364015.875p 0.552549mV 364016.428p 0.552549mV 364035.183p 0.55451mV 364051.097p 0.552142mV 364078.951p 0.5416mV 365003.576p 0.551981mV 365019.841p 0.552108mV 365021.806p 0.551663mV 365026.887p 0.550852mV 365106.666p 0.543638mV 365115.366p 0.542339mV 365117.762p 0.542339mV 365118.385p 0.542339mV 365123.638p 0.541137mV 366000.732p 0.55063mV 366016.118p 0.551845mV 366037.439p 0.554949mV 366068.479p 0.552009mV 366082.231p 0.546372mV 366115.347p 0.531156mV 367004.935p 0.550626mV 367006.152p 0.55062mV 367055.723p 0.555378mV 367058.574p 0.555378mV 367059.017p 0.555378mV 367065.067p 0.554307mV 367065.094p 0.554307mV 367100.042p 0.547885mV 367112.64p 0.545382mV 367116.455p 0.543948mV 368000.728p 0.547097mV 368017.787p 0.548426mV 368019.795p 0.548426mV 368062.117p 0.548811mV 368063.036p 0.548811mV 368070.814p 0.547896mV 368073.506p 0.547896mV 368076.607p 0.547988mV 368076.865p 0.547988mV 368077.111p 0.547988mV 368132.932p 0.552003mV 368145.201p 0.551258mV 369022.592p 0.54753mV 369038.334p 0.54397mV 370010.562p 0.554341mV 370016.502p 0.555134mV 370018.056p 0.555134mV 370027.18p 0.556358mV 370048.251p 0.558092mV 370049.581p 0.558092mV 370072.671p 0.552992mV 370078.282p 0.551611mV 370085.924p 0.547752mV 370103.127p 0.542141mV 371012.954p 0.554644mV 371013.876p 0.554644mV 371062.506p 0.557747mV 371065.762p 0.558544mV 371080.075p 0.562413mV 372029.072p 0.548874mV 372077.925p 0.546277mV 372078.105p 0.546277mV 372083.934p 0.547302mV 372097.047p 0.551849mV 372100.052p 0.553613mV 372104.358p 0.553613mV 373012.322p 0.547519mV 373022.624p 0.546246mV 373023.83p 0.546246mV 373034.921p 0.545705mV 373080.042p 0.537833mV 374012.279p 0.550805mV 374025.429p 0.549238mV 374054.893p 0.547071mV 374064.573p 0.54611mV 374110.865p 0.559299mV 374130.37p 0.568135mV 374131.101p 0.568135mV 374131.354p 0.568135mV 374133.283p 0.568135mV 374171.288p 0.590909mV 375020.671p 0.551738mV 375023.74p 0.551738mV 375030.608p 0.552759mV 376052.833p 0.545198mV 376071.151p 0.541882mV 376091.543p 0.540726mV 376103.207p 0.538669mV 377009.901p 0.548611mV 377013.323p 0.548991mV 377028.679p 0.550869mV 377046.903p 0.551691mV 377050.698p 0.552085mV 377053.461p 0.552085mV 377115.921p 0.536646mV 377134.231p 0.528787mV 378000.537p 0.547872mV 378017.043p 0.548804mV 378017.293p 0.548804mV 378021.847p 0.549116mV 378055.508p 0.552064mV 378060.4p 0.552389mV 378081.42p 0.550796mV 378086.445p 0.55004mV 378108.507p 0.544855mV 378111.403p 0.543747mV 378143.122p 0.539705mV 378170.562p 0.532084mV 378175.001p 0.529906mV 378184.689p 0.528096mV 378201.903p 0.518669mV 378236.982p 0.502312mV 378237.393p 0.502312mV 379039.004p 0.551434mV 379077.438p 0.554929mV 379121.12p 0.550231mV 379122.452p 0.550231mV 380016.944p 0.552695mV 380039.296p 0.553182mV 380093.68p 0.556826mV 380100.613p 0.557053mV 380128.61p 0.56109mV 380162.719p 0.567216mV 380166.107p 0.567891mV 380175.848p 0.568154mV 380239.976p 0.551681mV 380250.741p 0.549397mV 380261.987p 0.549692mV 380280.84p 0.549529mV 380288.566p 0.549484mV 380295.287p 0.550488mV 380347.731p 0.553267mV 380349.544p 0.553267mV 380352.306p 0.554313mV 381065.772p 0.555871mV 381074.84p 0.556192mV 382026.676p 0.54641mV 382027.094p 0.54641mV 382029.688p 0.54641mV 382032.694p 0.546037mV 382034.812p 0.546037mV 382036.779p 0.545297mV 382058.551p 0.54085mV 383024.812p 0.54528mV 383031.248p 0.543591mV 383049.19p 0.541243mV 384001.868p 0.551694mV 384038.488p 0.548348mV 384041.857p 0.546511mV 384049.078p 0.544306mV 385019.743p 0.54984mV 385019.799p 0.54984mV 385021.388p 0.551019mV 385044.554p 0.557199mV 386002.345p 0.551652mV 386014.319p 0.551328mV 386026.472p 0.55176mV 386029.997p 0.55176mV 386055.962p 0.553013mV 386061.673p 0.552677mV 386073.642p 0.550913mV 386086.947p 0.546993mV 386099.39p 0.545233mV 386112.22p 0.545329mV 387015.243p 0.553257mV 387017.267p 0.553257mV 387019.897p 0.553257mV 387031.102p 0.552359mV 387035.591p 0.551572mV 387077.464p 0.542293mV 388004.367p 0.547914mV 388023.904p 0.547581mV 388030.817p 0.546316mV 388047.564p 0.5435mV 388072.864p 0.541948mV 388126.973p 0.541796mV 388137.005p 0.543349mV 388140.313p 0.543572mV 389011.651p 0.553973mV 389034.751p 0.556556mV 389034.903p 0.556556mV 389045.317p 0.558879mV 389062.463p 0.558673mV 390011.026p 0.551204mV 390014.204p 0.551204mV 390016.586p 0.551162mV 390023.109p 0.551485mV 390030.482p 0.551766mV 390043.13p 0.552046mV 390083.988p 0.563432mV 391002.975p 0.546561mV 391077.946p 0.536217mV 392009.511p 0.553492mV 392013.081p 0.553837mV 392015.6p 0.554548mV 392017.546p 0.554548mV 392032.739p 0.556683mV 392040.106p 0.557013mV 392042.644p 0.557013mV 392043.42p 0.557013mV 393003.002p 0.55176mV 393010.012p 0.552222mV 393025.381p 0.554921mV 393029.438p 0.554921mV 393060.713p 0.558906mV 394017.121p 0.545589mV 394046.53p 0.546998mV 394099.87p 0.549772mV 396017.536p 0.554254mV 396023.063p 0.55388mV 396031.409p 0.552762mV 396050.146p 0.55124mV 397001.866p 0.554527mV 397038.67p 0.556404mV 398033.087p 0.545973mV 398077.703p 0.546597mV 398083.595p 0.546293mV 399008.597p 0.550518mV 399036.381p 0.552747mV 399045.934p 0.554471mV 399060.806p 0.556521mV 399068.135p 0.557209mV 400024.541p 0.54503mV 400029.238p 0.545051mV 400045.852p 0.546578mV 400073.021p 0.549915mV 400082.375p 0.551023mV 400084.219p 0.551023mV 400084.568p 0.551023mV 400100.252p 0.556158mV 400121.726p 0.563494mV 400130.746p 0.566079mV 401067.246p 0.556147mV 401074.559p 0.556491mV 401079.922p 0.556472mV 401101.303p 0.553874mV 401118.499p 0.551333mV 401128.945p 0.550263mV 401145.648p 0.547426mV 401166.567p 0.546832mV 401168.102p 0.546832mV 401172.564p 0.54724mV 402074.772p 0.552674mV 402077.436p 0.552715mV 402079.212p 0.552715mV 402083.873p 0.55312mV 402098.229p 0.554324mV 402126.228p 0.554855mV 402139.666p 0.555988mV 402168.936p 0.560062mV 402172.936p 0.560427mV 402178.791p 0.560425mV 402179.247p 0.560425mV 402180.952p 0.560056mV 403043.897p 0.549159mV 403051.603p 0.550224mV 403061.102p 0.550562mV 403084.254p 0.549789mV 403105.454p 0.544633mV 403133.925p 0.544217mV 403157.021p 0.543401mV 403192.604p 0.54028mV 403196.36p 0.54024mV 403210.108p 0.539366mV 404042.979p 0.543354mV 404045.4p 0.542603mV 404046.49p 0.542603mV 405014.666p 0.546095mV 405051.061p 0.54759mV 405060.067p 0.550153mV 405080.004p 0.555286mV 406006.242p 0.547716mV 406008.891p 0.547716mV 406011.414p 0.547366mV 406030.667p 0.545222mV 406037.297p 0.544499mV 406071.849p 0.544479mV 406084.012p 0.545539mV 406098.981p 0.548751mV 406109.898p 0.551974mV 406142.894p 0.561196mV 406204.055p 0.575368mV 406231.497p 0.583657mV 407022.919p 0.550224mV 407037.994p 0.548317mV 407044.458p 0.547194mV 407051.388p 0.544581mV 407055.767p 0.543822mV 407056.841p 0.543822mV 407057.511p 0.543822mV 407079.706p 0.540767mV 407080.0p 0.540767mV 407095.755p 0.538402mV 408044.161p 0.551616mV 408062.23p 0.550276mV 408071.43p 0.549238mV 408081.943p 0.54893mV 408110.612p 0.550178mV 408146.112p 0.554345mV 408147.288p 0.554345mV 408170.034p 0.558476mV 409023.588p 0.547056mV 409038.168p 0.541823mV 410006.546p 0.552267mV 410008.91p 0.552267mV 410016.572p 0.553196mV 410031.074p 0.555864mV 410044.969p 0.557521mV 411013.732p 0.553406mV 412005.447p 0.554157mV 412013.573p 0.553729mV 412037.856p 0.552699mV 412070.889p 0.554519mV 413000.541p 0.549114mV 413000.842p 0.549114mV 413008.454p 0.549198mV 413033.73p 0.550735mV 413047.377p 0.54846mV 413057.718p 0.546829mV 413059.284p 0.546829mV 413117.665p 0.550265mV 413140.087p 0.545386mV 413168.615p 0.538744mV 413177.135p 0.535729mV 413181.607p 0.53404mV 413190.128p 0.531759mV 413190.212p 0.531759mV 413195.012p 0.530435mV 413204.873p 0.528745mV 413208.662p 0.52742mV 414055.541p 0.547725mV 414060.598p 0.548859mV 414077.585p 0.55079mV 414089.064p 0.553413mV 414104.083p 0.557162mV 414139.789p 0.564364mV 414160.81p 0.566447mV 414184.921p 0.566711mV 414190.412p 0.568692mV 414198.276p 0.570235mV 415030.046p 0.551989mV 415041.632p 0.556715mV 416004.304p 0.551888mV 416006.589p 0.551965mV 416029.309p 0.550064mV 416035.126p 0.54764mV 416055.834p 0.545682mV 416066.335p 0.546869mV 416069.994p 0.546869mV 416074.701p 0.547274mV 416079.604p 0.547309mV 417047.897p 0.546008mV 417048.129p 0.546008mV 418041.28p 0.54913mV 418053.229p 0.549417mV 419006.245p 0.552249mV 419023.651p 0.551395mV 420031.235p 0.547968mV 420049.024p 0.547672mV 420069.284p 0.549949mV 420095.587p 0.553361mV 420100.902p 0.55448mV 420126.814p 0.561929mV 421008.995p 0.545242mV 421012.427p 0.544791mV 421065.309p 0.53827mV 421081.645p 0.53793mV 421082.32p 0.53793mV 421089.335p 0.537808mV 422008.789p 0.547547mV 422055.044p 0.552958mV 422073.439p 0.557138mV 423005.296p 0.545997mV 423010.401p 0.546357mV 423014.414p 0.546357mV 423021.246p 0.547446mV 423040.262p 0.548182mV 423042.931p 0.548182mV 423093.957p 0.54361mV 423127.052p 0.537647mV 423133.94p 0.537321mV 423138.517p 0.53663mV 423138.677p 0.53663mV 423163.431p 0.535014mV 423168.679p 0.535791mV 423172.54p 0.536935mV 423174.317p 0.536935mV 423188.506p 0.539648mV 424000.149p 0.546171mV 424001.839p 0.546171mV 424005.107p 0.54625mV 424009.643p 0.54625mV 424019.269p 0.545308mV 424028.279p 0.542898mV 424032.52p 0.541142mV 424044.5p 0.537989mV 425032.567p 0.552683mV 425035.6p 0.553489mV 425035.936p 0.553489mV 425053.075p 0.553727mV 425053.543p 0.553727mV 425101.254p 0.545504mV 425151.551p 0.539494mV 425151.74p 0.539494mV 425164.429p 0.536385mV 426054.017p 0.54525mV 427050.726p 0.543675mV 428005.02p 0.548576mV 428019.923p 0.549552mV 428021.278p 0.549857mV 428022.155p 0.549857mV 428026.43p 0.549797mV 428114.146p 0.53602mV 429002.825p 0.545807mV 429011.595p 0.545614mV 429020.352p 0.544691mV 429039.259p 0.54532mV 429067.098p 0.549143mV 429090.183p 0.558029mV 429094.317p 0.558029mV 430010.104p 0.547043mV 430018.422p 0.546286mV 430027.888p 0.543674mV 430032.957p 0.541817mV 430037.58p 0.539594mV 431037.597p 0.542433mV 431072.314p 0.548811mV 431081.447p 0.550591mV 431094.498p 0.55165mV 431099.727p 0.552367mV 432004.737p 0.548618mV 432026.689p 0.546819mV 432031.11p 0.546382mV 432031.596p 0.546382mV 432055.787p 0.543074mV 432060.817p 0.541893mV 433001.293p 0.5489mV 433016.27p 0.550153mV 433022.395p 0.550573mV 433053.185p 0.553502mV 434003.679p 0.546675mV 434006.525p 0.546644mV 434011.112p 0.54698mV 434016.326p 0.547682mV 434035.418p 0.55416mV 435000.016p 0.553189mV 436031.722p 0.552564mV 436032.827p 0.552564mV 436079.598p 0.553857mV 436080.071p 0.552832mV 436097.936p 0.547574mV 437008.76p 0.552016mV 437012.45p 0.551722mV 437027.745p 0.55303mV 437034.202p 0.554197mV 437036.925p 0.555729mV 437041.03p 0.556896mV 437046.713p 0.558429mV 437067.054p 0.563844mV 438002.34p 0.553075mV 438014.209p 0.553506mV 438015.446p 0.55354mV 438026.688p 0.553247mV 438028.936p 0.553247mV 438040.736p 0.551903mV 438068.465p 0.554318mV 438075.238p 0.554782mV 438090.687p 0.556411mV 439011.283p 0.548617mV 439013.433p 0.548617mV 439020.177p 0.548354mV 439081.348p 0.544581mV 439087.414p 0.544629mV 439097.972p 0.544354mV 439126.722p 0.544948mV 439161.88p 0.553177mV 439164.108p 0.553177mV 439172.465p 0.557977mV 439181.434p 0.563513mV 439182.803p 0.563513mV 439186.636p 0.565737mV 440090.477p 0.558556mV 441043.525p 0.545935mV 441053.554p 0.542672mV 442049.312p 0.543737mV 443000.579p 0.551864mV 443004.317p 0.551864mV 443026.901p 0.552534mV 443082.105p 0.561075mV 443086.462p 0.561784mV 444000.605p 0.553118mV 444003.323p 0.553118mV 444035.537p 0.551863mV 444062.43p 0.546299mV 444071.913p 0.54371mV 444108.937p 0.541001mV 444115.112p 0.542036mV 444162.58p 0.554493mV 445011.126p 0.550117mV 445033.771p 0.552221mV 445047.168p 0.555447mV 445069.639p 0.55977mV 445073.085p 0.561588mV 446033.521p 0.556113mV 446034.968p 0.556113mV 446035.571p 0.557492mV 447000.899p 0.547413mV 447014.045p 0.547155mV 447022.572p 0.545432mV 447027.722p 0.54402mV 448059.855p 0.560557mV 449033.982p 0.54798mV 449034.614p 0.54798mV 449073.413p 0.552992mV 449073.909p 0.552992mV 449078.389p 0.55453mV 449133.069p 0.562766mV 449137.143p 0.563597mV 450011.57p 0.546492mV 450012.313p 0.546492mV 450012.495p 0.546492mV 450015.35p 0.546484mV 450041.814p 0.540936mV 451017.273p 0.55505mV 451041.944p 0.555025mV 451066.482p 0.561971mV 451071.013p 0.563731mV 452006.103p 0.549211mV 452028.643p 0.549916mV 452075.776p 0.545158mV 452113.798p 0.537839mV 452118.741p 0.53637mV 453005.867p 0.547706mV 453019.001p 0.547413mV 453020.604p 0.547082mV 453031.194p 0.547513mV 453034.863p 0.547513mV 453074.128p 0.553589mV 453086.411p 0.554772mV 453089.96p 0.554772mV 453117.915p 0.553861mV 453121.662p 0.553528mV 453148.146p 0.555149mV 453169.948p 0.560396mV 453177.977p 0.564489mV 454032.202p 0.557115mV 455002.636p 0.55425mV 455019.267p 0.554454mV 455050.388p 0.554117mV 455065.129p 0.557284mV 455065.92p 0.557284mV 455089.869p 0.561542mV 456002.067p 0.553734mV 456003.53p 0.553734mV 456016.556p 0.555038mV 456024.756p 0.556203mV 456034.856p 0.557437mV 457024.726p 0.554095mV 457032.768p 0.556488mV 457042.888p 0.558157mV 458014.484p 0.554319mV 458021.915p 0.553238mV 459008.73p 0.549283mV 459043.532p 0.553987mV 459055.784p 0.55786mV 460022.0p 0.544306mV 460025.802p 0.542924mV 460026.373p 0.542924mV 460047.027p 0.538855mV 461000.191p 0.552578mV 461008.143p 0.552543mV 461022.127p 0.55243mV 462003.763p 0.546277mV 462015.265p 0.54644mV 462030.577p 0.546242mV 462065.518p 0.554225mV 463004.469p 0.553874mV 463012.828p 0.554191mV 463050.04p 0.562792mV 464032.238p 0.552007mV 464069.772p 0.556373mV 464085.389p 0.559138mV 465007.788p 0.551351mV 465021.016p 0.552598mV 465031.908p 0.554285mV 465036.037p 0.554946mV 466014.372p 0.550921mV 466036.324p 0.554838mV 466052.055p 0.559404mV 467025.545p 0.550281mV 468023.381p 0.546299mV 468045.612p 0.554019mV 468053.831p 0.55593mV 468056.174p 0.557479mV 468059.584p 0.557479mV 468061.346p 0.558664mV 469037.472p 0.54045mV 469037.503p 0.54045mV 469066.302p 0.53226mV 470018.12p 0.551934mV 470029.632p 0.551566mV 470040.576p 0.551556mV 470045.009p 0.551552mV 470051.831p 0.551181mV 470083.058p 0.555151mV 470094.139p 0.55696mV 470105.522p 0.560958mV 470111.676p 0.562051mV 470119.288p 0.56278mV 470126.76p 0.564613mV 470127.092p 0.564613mV 470131.896p 0.565718mV 471000.955p 0.554269mV 471008.045p 0.554324mV 471017.324p 0.554802mV 471023.046p 0.555225mV 471043.353p 0.556929mV 471046.176p 0.557724mV 471067.393p 0.563849mV 472054.034p 0.539431mV 473003.433p 0.545358mV 473043.387p 0.543155mV 473061.678p 0.540185mV 473072.967p 0.538318mV 474023.06p 0.547018mV 474035.626p 0.550104mV 474036.974p 0.550104mV 475020.835p 0.547866mV 475040.228p 0.545727mV 475061.959p 0.544297mV 475062.558p 0.544297mV 476022.032p 0.548182mV 476047.889p 0.546368mV 476049.902p 0.546368mV 476050.158p 0.54593mV 476074.132p 0.545626mV 477010.298p 0.549624mV 477062.654p 0.541343mV 477073.002p 0.538639mV 478015.77p 0.547839mV 478039.362p 0.546961mV 478094.246p 0.554561mV 478097.614p 0.555986mV 478113.642p 0.561739mV 478114.704p 0.561739mV 479045.252p 0.545239mV 479060.841p 0.547226mV 479066.398p 0.547892mV 480001.402p 0.550528mV 480014.703p 0.550187mV 480068.645p 0.556588mV 481003.956p 0.547075mV 481009.14p 0.547097mV 481020.001p 0.546425mV 481055.585p 0.551276mV 481064.362p 0.553116mV 481067.297p 0.554591mV 481083.417p 0.558292mV 481092.765p 0.561624mV 481093.144p 0.561624mV 482013.067p 0.552325mV 482018.729p 0.551558mV 482071.551p 0.538752mV 483008.737p 0.545747mV 483024.348p 0.545782mV 483044.031p 0.542891mV 484004.429p 0.545343mV 484008.514p 0.545413mV 484057.116p 0.544235mV 484080.029p 0.545595mV 484088.824p 0.545642mV 484092.905p 0.546051mV 484112.11p 0.546203mV 484129.791p 0.546653mV 484141.235p 0.548165mV 484150.037p 0.549275mV 484159.875p 0.550005mV 484161.057p 0.551096mV 484171.305p 0.552899mV 484177.009p 0.55361mV 485009.759p 0.552854mV 485043.587p 0.554302mV 485077.865p 0.553169mV 485101.372p 0.552761mV 485110.316p 0.553105mV 485111.789p 0.553105mV 485143.125p 0.559232mV 485150.2p 0.563224mV 485167.436p 0.568678mV 485169.102p 0.568678mV 486034.446p 0.548613mV 487019.114p 0.546042mV 487043.474p 0.540371mV 487050.555p 0.537722mV 487052.765p 0.537722mV 488007.12p 0.546499mV 488019.848p 0.545971mV 488079.589p 0.552331mV 488093.085p 0.55432mV 488094.007p 0.55432mV 489013.697p 0.546854mV 489016.771p 0.546787mV 489019.863p 0.546787mV 489067.437p 0.54502mV 489075.791p 0.544519mV 489091.074p 0.545775mV 489126.514p 0.544178mV 489184.74p 0.541841mV 489208.846p 0.539902mV 489208.965p 0.539902mV 489211.123p 0.539432mV 490021.274p 0.554025mV 490026.07p 0.554723mV 490041.0p 0.556087mV 490064.694p 0.55669mV 490096.284p 0.553202mV 490121.932p 0.542456mV 491018.436p 0.553349mV 492053.062p 0.557188mV 492056.414p 0.557972mV 492064.175p 0.558395mV 493018.671p 0.547832mV 493056.557p 0.542003mV 494016.428p 0.547173mV 494042.393p 0.547235mV 495001.854p 0.550602mV 495064.191p 0.551489mV 495070.012p 0.551053mV 495085.571p 0.548404mV 495099.652p 0.546527mV 495100.441p 0.545407mV 495104.981p 0.545407mV 495108.42p 0.544655mV 495128.299p 0.545313mV 496006.131p 0.553411mV 496015.422p 0.553655mV 496055.618p 0.561189mV 497056.508p 0.549491mV 497057.35p 0.549491mV 497069.107p 0.55054mV 497072.759p 0.550886mV 497083.735p 0.550487mV 497091.074p 0.550831mV 497118.422p 0.550105mV 497138.801p 0.546526mV 497143.821p 0.545459mV 497222.576p 0.516359mV 497250.798p 0.504689mV 497291.735p 0.488309mV 498040.711p 0.557944mV 498057.465p 0.556811mV 498058.461p 0.556811mV 498076.117p 0.553146mV 498081.46p 0.552784mV 499021.629p 0.554453mV 499025.416p 0.555915mV 500002.427p 0.55011mV 500007.242p 0.550124mV 500029.942p 0.547979mV 500030.923p 0.546891mV 500032.66p 0.546891mV 500036.293p 0.546167mV 500053.18p 0.542521mV 500053.664p 0.542521mV 502003.763p 0.55071mV 502018.627p 0.551056mV 502034.712p 0.549568mV 502057.793p 0.550245mV 502066.512p 0.550583mV 502081.037p 0.548342mV 502082.4p 0.548342mV 502091.904p 0.547209mV 502092.876p 0.547209mV 502110.896p 0.545649mV 502124.62p 0.545218mV 502140.766p 0.546506mV 502144.146p 0.546506mV 502151.309p 0.546763mV 502158.999p 0.546703mV 502173.337p 0.547956mV 502175.238p 0.547878mV 502176.935p 0.547878mV 503016.542p 0.553897mV 504000.058p 0.549623mV 504007.664p 0.549639mV 504013.364p 0.549289mV 504021.204p 0.549684mV 504027.1p 0.549698mV 504052.187p 0.550124mV 504066.404p 0.551248mV 504073.229p 0.552353mV 504076.179p 0.553092mV 504089.749p 0.555668mV 504090.567p 0.556774mV 504093.817p 0.556774mV 505003.337p 0.550428mV 505014.55p 0.550813mV 505033.127p 0.555974mV 505033.979p 0.555974mV 505044.555p 0.560023mV 506008.193p 0.552303mV 506029.931p 0.552603mV 506039.402p 0.553848mV 506042.223p 0.55502mV 506053.957p 0.55773mV 506072.877p 0.559511mV 506102.511p 0.564824mV 507028.227p 0.551031mV 508008.054p 0.551329mV 508019.252p 0.550206mV 508022.585p 0.549097mV 508048.125p 0.540254mV 508051.77p 0.538407mV 509014.875p 0.551967mV 509034.434p 0.554276mV 509035.158p 0.554305mV 509035.36p 0.554305mV 509046.274p 0.553265mV 509060.808p 0.548963mV 509070.477p 0.544993mV 509074.017p 0.544993mV 510004.643p 0.553731mV 510025.362p 0.55377mV 510052.727p 0.552009mV 510087.498p 0.547378mV 510094.92p 0.547029mV 510134.342p 0.550055mV 510134.813p 0.550055mV 510156.672p 0.548651mV 510164.188p 0.548298mV 510168.687p 0.54758mV 510204.973p 0.546929mV 510246.221p 0.554331mV 510247.858p 0.554331mV 511015.729p 0.547805mV 511026.195p 0.546878mV 511033.344p 0.546599mV 511056.543p 0.54338mV 511060.073p 0.54237mV 511065.368p 0.540994mV 511077.991p 0.537871mV 511094.769p 0.532985mV 511094.786p 0.532985mV 512041.465p 0.555355mV 512130.285p 0.557482mV 512132.363p 0.557482mV 512189.693p 0.539191mV 512201.358p 0.532762mV 512252.917p 0.520537mV 512264.616p 0.517374mV 512265.301p 0.515247mV 512301.162p 0.494545mV 513002.096p 0.552958mV 513031.367p 0.550817mV 513074.589p 0.543995mV 514015.056p 0.555317mV 514020.511p 0.556374mV 514041.248p 0.562075mV 514062.171p 0.566352mV 515003.872p 0.546789mV 515025.08p 0.542785mV 515032.715p 0.541619mV 515041.146p 0.538919mV 515041.36p 0.538919mV 515049.318p 0.538116mV 515074.05p 0.532228mV 516002.358p 0.554671mV 516014.735p 0.555097mV 516055.388p 0.559096mV 516079.091p 0.560777mV 516089.84p 0.559813mV 516093.35p 0.55952mV 516129.499p 0.555403mV 516135.219p 0.552342mV 516136.616p 0.552342mV 516137.98p 0.552342mV 516143.008p 0.550635mV 516146.457p 0.548569mV 516178.108p 0.541001mV 517034.473p 0.544323mV 517040.558p 0.542499mV 518016.983p 0.544992mV 518026.48p 0.543106mV 518059.177p 0.535214mV 519032.562p 0.551956mV 519052.512p 0.555204mV 519072.45p 0.557733mV 519089.804p 0.557635mV 519091.697p 0.557362mV 520010.14p 0.54787mV 520013.411p 0.54787mV 520028.183p 0.548934mV 520050.91p 0.548534mV 520076.22p 0.549265mV 520112.997p 0.549355mV 520128.819p 0.549805mV 521024.817p 0.549306mV 521047.223p 0.551549mV 521072.834p 0.557115mV 521079.913p 0.558601mV 521080.931p 0.559725mV 522004.457p 0.553252mV 522005.42p 0.553332mV 522033.295p 0.557749mV 522040.111p 0.559736mV 522045.444p 0.561279mV 522072.143p 0.567939mV 523012.487p 0.549212mV 523030.843p 0.552328mV 523075.625p 0.55575mV 524012.579p 0.553335mV 524029.272p 0.550206mV 525015.025p 0.554122mV 525038.152p 0.551203mV 525040.898p 0.550105mV 525063.707p 0.542773mV 526063.642p 0.553021mV 526092.816p 0.556833mV 526094.629p 0.556833mV 526116.435p 0.560332mV 526120.241p 0.561402mV 527019.163p 0.547166mV 527022.257p 0.546125mV 527038.383p 0.540808mV 527046.055p 0.536892mV 527049.089p 0.536892mV 528002.052p 0.551078mV 528085.037p 0.549752mV 528092.704p 0.550158mV 528128.477p 0.555132mV 528134.643p 0.556254mV 528163.484p 0.566997mV 528183.785p 0.572968mV 529032.871p 0.551367mV 529042.513p 0.54942mV 530002.493p 0.554643mV 530006.703p 0.554554mV 530026.279p 0.552726mV 530035.638p 0.551438mV 530047.407p 0.54868mV 531037.121p 0.554157mV 531046.847p 0.554672mV 531081.525p 0.551546mV 531083.324p 0.551546mV 531110.828p 0.545027mV 532011.459p 0.551097mV 532051.497p 0.556322mV 532057.205p 0.556984mV 532133.77p 0.544017mV 532138.695p 0.541819mV 532161.075p 0.530501mV 532174.422p 0.525765mV 533011.228p 0.548111mV 533023.31p 0.549047mV 533077.375p 0.550735mV 534006.277p 0.550114mV 534014.657p 0.549678mV 534017.821p 0.548877mV 534021.3p 0.548443mV 534038.074p 0.54568mV 534056.952p 0.538822mV 535004.725p 0.548026mV 535015.699p 0.54824mV 535023.47p 0.548555mV 535076.477p 0.549857mV 535099.857p 0.546767mV 535105.123p 0.544862mV 535113.256p 0.543727mV 535115.776p 0.542958mV 535148.834p 0.532835mV 535150.098p 0.530227mV 536028.577p 0.549004mV 536044.914p 0.549653mV 536049.721p 0.550358mV 536073.731p 0.5506mV 536075.916p 0.550579mV 536086.308p 0.550905mV 536102.649p 0.552316mV 536108.749p 0.552302mV 536122.964p 0.554467mV 536131.59p 0.557749mV 537029.915p 0.550179mV 537038.11p 0.550432mV 537055.066p 0.551674mV 537056.144p 0.551674mV 537064.726p 0.551254mV 537068.526p 0.551202mV 537074.154p 0.551516mV 538019.801p 0.548368mV 538023.571p 0.54873mV 538057.382p 0.55272mV 538059.205p 0.55272mV 538062.242p 0.553814mV 539037.959p 0.550179mV 539047.154p 0.551372mV 539055.371p 0.553302mV 540016.262p 0.55371mV 540033.205p 0.551251mV 540034.503p 0.551251mV 540076.405p 0.548302mV 540104.108p 0.546802mV 540116.106p 0.546202mV 540153.446p 0.549347mV 540155.1p 0.550013mV 541020.417p 0.554301mV 541030.732p 0.554777mV 541039.999p 0.554834mV 541062.202p 0.557699mV 541071.389p 0.558202mV 541073.121p 0.558202mV 541078.562p 0.559005mV 541082.795p 0.559446mV 541103.825p 0.559785mV 542047.136p 0.55457mV 542066.478p 0.554077mV 542066.969p 0.554077mV 543006.933p 0.550949mV 543021.791p 0.550782mV 543026.59p 0.550728mV 543029.723p 0.550728mV 543036.295p 0.550256mV 543039.931p 0.550256mV 543040.025p 0.549838mV 543046.565p 0.549055mV 543158.524p 0.54353mV 543181.062p 0.555061mV 544006.216p 0.547645mV 544012.533p 0.547997mV 544027.775p 0.548329mV 544029.997p 0.548329mV 544037.157p 0.547215mV 544071.761p 0.547925mV 544108.115p 0.547611mV 544111.082p 0.547993mV 545002.684p 0.550493mV 545006.317p 0.550484mV 545006.442p 0.550484mV 545029.687p 0.551182mV 545030.997p 0.55154mV 545095.152p 0.55225mV 545097.482p 0.55225mV 545108.806p 0.554824mV 545119.584p 0.556676mV 546025.305p 0.545756mV 547039.973p 0.546936mV 547055.795p 0.540377mV 547063.53p 0.537819mV 548018.22p 0.549125mV 548049.828p 0.554189mV 548079.834p 0.551956mV 548091.566p 0.550666mV 549008.401p 0.54541mV 549015.571p 0.545634mV 549018.445p 0.545634mV 549040.784p 0.54417mV 549044.562p 0.54417mV 549090.169p 0.550316mV 550044.112p 0.550585mV 550052.641p 0.547462mV 550057.885p 0.54535mV 551015.471p 0.553603mV 551016.759p 0.553603mV 551030.367p 0.551909mV 552053.524p 0.546123mV 552054.08p 0.546123mV 552059.989p 0.544619mV 552069.558p 0.541238mV 553016.82p 0.547902mV 553040.627p 0.547867mV 553066.922p 0.54967mV 553067.271p 0.54967mV 553071.008p 0.550106mV 553095.061p 0.557793mV 554000.891p 0.548154mV 554005.75p 0.548213mV 554033.299p 0.553988mV 555020.876p 0.544911mV 555023.671p 0.544911mV 555028.135p 0.544154mV 555029.053p 0.544154mV 556009.048p 0.550988mV 556017.727p 0.550709mV 556045.403p 0.549146mV 556049.743p 0.549146mV 556064.958p 0.544887mV 557008.477p 0.548735mV 557013.957p 0.548382mV 557036.044p 0.546987mV 557053.752p 0.546298mV 557061.29p 0.544496mV 557070.025p 0.541228mV 558011.174p 0.549003mV 558011.588p 0.549003mV 558018.181p 0.548351mV 558060.115p 0.54285mV 559015.475p 0.549787mV 559032.662p 0.549684mV 559068.253p 0.549794mV 559095.153p 0.555046mV 559096.435p 0.555046mV 559127.161p 0.563262mV 560013.127p 0.551821mV 560013.575p 0.551821mV 560019.615p 0.55107mV 560025.044p 0.549206mV 560031.113p 0.548823mV 560057.363p 0.542877mV 561026.307p 0.547883mV 561030.07p 0.546849mV 561030.95p 0.546849mV 561043.795p 0.544413mV 562018.835p 0.545588mV 562050.894p 0.540922mV 562051.174p 0.540922mV 562099.587p 0.5281mV 563018.02p 0.551129mV 563034.962p 0.549941mV 563063.823p 0.550858mV 563088.721p 0.554978mV 563102.262p 0.559658mV 564005.382p 0.550309mV 564015.621p 0.550683mV 564061.645p 0.544481mV 564070.055p 0.542641mV 565031.337p 0.557768mV 566000.449p 0.547529mV 566027.463p 0.543463mV 566038.232p 0.540011mV 566052.201p 0.536105mV 567019.457p 0.54778mV 567033.309p 0.548251mV 567105.731p 0.555332mV 567116.266p 0.555541mV 567116.437p 0.555541mV 567126.597p 0.554296mV 567170.705p 0.548954mV 567181.506p 0.549201mV 567181.735p 0.549201mV 567187.561p 0.549875mV 567199.223p 0.551591mV 567209.536p 0.553316mV 567218.919p 0.555052mV 568007.201p 0.55245mV 568030.426p 0.551549mV 568053.38p 0.548031mV 568057.049p 0.546598mV 568059.697p 0.546598mV 569000.606p 0.551858mV 569016.9p 0.550716mV 569038.587p 0.54699mV 569042.756p 0.545873mV 569043.639p 0.545873mV 570067.364p 0.560486mV 571023.834p 0.547932mV 571028.257p 0.547988mV 571043.354p 0.549623mV 571057.534p 0.553099mV 572010.021p 0.548546mV 572018.918p 0.547733mV 572043.542p 0.54697mV 572045.823p 0.546892mV 572062.375p 0.548853mV 572065.873p 0.55024mV 573018.864p 0.551822mV 574043.012p 0.551674mV 574086.973p 0.548339mV 574093.528p 0.548013mV 574102.232p 0.546995mV 574107.998p 0.546303mV 574119.396p 0.543821mV 574132.034p 0.540272mV 574134.011p 0.540272mV 574135.888p 0.538841mV 574136.606p 0.538841mV 574137.744p 0.538841mV 575015.95p 0.549636mV 575026.58p 0.550912mV 575027.587p 0.550912mV 575042.574p 0.555581mV 576007.73p 0.547495mV 576041.022p 0.548261mV 576078.374p 0.550872mV 576080.19p 0.551251mV 576123.82p 0.548508mV 576130.725p 0.547478mV 576136.374p 0.546782mV 576156.896p 0.541821mV 576160.069p 0.540765mV 576170.553p 0.539753mV 576192.083p 0.536998mV 576214.464p 0.53278mV 576227.398p 0.528877mV 577021.569p 0.550891mV 577046.472p 0.547667mV 577057.655p 0.547461mV 577069.683p 0.547245mV 577101.704p 0.549128mV 577139.733p 0.55411mV 577158.242p 0.557066mV 578020.854p 0.552337mV 578031.921p 0.552571mV 578060.227p 0.548857mV 579056.695p 0.550482mV 579071.36p 0.546015mV 580055.651p 0.551373mV 580061.3p 0.549595mV 580092.892p 0.546573mV 580124.839p 0.55004mV 580145.868p 0.550127mV 580170.78p 0.548329mV 580175.976p 0.548324mV 580185.16p 0.548666mV 580188.452p 0.548666mV 581013.73p 0.552255mV 581027.586p 0.550923mV 581033.706p 0.550478mV 581045.805p 0.548408mV 581051.519p 0.54796mV 581055.846p 0.547145mV 581082.84p 0.543408mV 582005.36p 0.548841mV 582013.635p 0.548426mV 582023.361p 0.546496mV 582056.517p 0.54424mV 582059.611p 0.54424mV 582073.657p 0.541814mV 583016.561p 0.547056mV 583024.486p 0.546718mV 583048.327p 0.541018mV 583057.701p 0.538516mV 584008.271p 0.546728mV 584016.534p 0.546261mV 584061.683p 0.545378mV 584063.031p 0.545378mV 585018.119p 0.554811mV 585023.42p 0.555929mV 585037.609p 0.558554mV 585044.495p 0.559677mV 585051.344p 0.560832mV 587019.072p 0.548808mV 587043.388p 0.54842mV 587064.251p 0.549142mV 587120.864p 0.552895mV 587159.422p 0.550573mV 589010.646p 0.553035mV 589015.262p 0.553023mV 589033.627p 0.552992mV 589046.691p 0.556261mV 589074.24p 0.561754mV 589078.595p 0.56177mV 590027.528p 0.549447mV 590044.024p 0.553855mV 590049.157p 0.555328mV 591015.886p 0.551125mV 591042.588p 0.550271mV 591052.233p 0.551465mV 591059.901p 0.551514mV 591080.907p 0.551399mV 591101.996p 0.551608mV 591108.264p 0.551661mV 591125.461p 0.551883mV 591154.203p 0.554011mV 591156.416p 0.555538mV 591161.147p 0.557432mV 592002.989p 0.552456mV 592026.402p 0.553939mV 592047.607p 0.559812mV 592056.717p 0.561661mV 592066.732p 0.562791mV 592074.019p 0.56391mV 592084.984p 0.565064mV 593021.207p 0.551541mV 594001.356p 0.550391mV 594005.217p 0.550332mV 594014.309p 0.549907mV 594062.846p 0.544486mV 595010.002p 0.5487mV 595034.995p 0.549615mV 595087.109p 0.558518mV 595096.931p 0.559723mV 595107.554p 0.56167mV 596007.804p 0.547678mV 596039.046p 0.546997mV 596059.715p 0.545781mV 596075.622p 0.543794mV 597002.375p 0.549186mV 597010.539p 0.548823mV 597012.367p 0.548823mV 597029.457p 0.547739mV 597068.296p 0.544146mV 597081.063p 0.542708mV 597090.407p 0.543089mV 597103.636p 0.542736mV 597125.43p 0.545691mV 597134.759p 0.546795mV 597135.335p 0.547534mV 597138.017p 0.547534mV 597140.837p 0.547909mV 597188.717p 0.548112mV 598037.677p 0.549184mV 599018.734p 0.552776mV 599030.871p 0.554752mV 599071.839p 0.550575mV 600062.255p 0.56185mV 601070.207p 0.549574mV 601158.745p 0.568407mV 602013.738p 0.552598mV 602027.191p 0.549227mV 602034.416p 0.548103mV 602035.698p 0.547342mV 602039.303p 0.547342mV 602051.32p 0.544317mV 602061.593p 0.541676mV 603051.809p 0.543717mV 604012.26p 0.546477mV 604022.667p 0.546906mV 604036.766p 0.549569mV 604051.966p 0.553348mV 605009.581p 0.549491mV 605028.361p 0.552064mV 605084.49p 0.547441mV 605110.592p 0.547248mV 605114.633p 0.547248mV 605125.905p 0.55024mV 605136.447p 0.55406mV 605143.762p 0.55652mV 605145.802p 0.559346mV 606014.19p 0.552174mV 606015.165p 0.552125mV 606035.636p 0.553392mV 606057.562p 0.549542mV 606065.336p 0.547616mV 606084.197p 0.545996mV 606105.53p 0.545687mV 606122.844p 0.546197mV 606135.235p 0.547047mV 606147.128p 0.545771mV 606163.005p 0.544745mV 607000.31p 0.549538mV 607001.398p 0.549538mV 607012.195p 0.549848mV 607015.798p 0.550552mV 607022.277p 0.551621mV 607041.602p 0.559564mV 608006.796p 0.551899mV 608012.071p 0.551517mV 608085.995p 0.540579mV 608101.477p 0.542617mV 608102.416p 0.542617mV 608116.24p 0.54571mV 608136.005p 0.546856mV 608139.053p 0.546856mV 609040.1p 0.549543mV 610027.035p 0.551943mV 610052.135p 0.55477mV 610076.148p 0.556497mV 610091.872p 0.558421mV 610092.039p 0.558421mV 610101.303p 0.559344mV 610110.092p 0.561006mV 611008.928p 0.550812mV 611011.693p 0.551194mV 611045.061p 0.556798mV 612009.924p 0.552143mV 613005.185p 0.553609mV 613032.74p 0.54955mV 613064.839p 0.544704mV 614032.349p 0.546867mV 614053.968p 0.543318mV 615013.068p 0.545516mV 615025.85p 0.543198mV 615028.676p 0.543198mV 615055.124p 0.539634mV 616031.702p 0.551345mV 616042.792p 0.551598mV 616082.508p 0.548999mV 616083.302p 0.548999mV 616092.343p 0.545619mV 616098.791p 0.543381mV 616108.241p 0.540001mV 617030.594p 0.545489mV 617062.738p 0.545977mV 617073.585p 0.544181mV 617099.004p 0.539106mV 618003.103p 0.554373mV 618044.792p 0.553289mV 618045.097p 0.553248mV 618079.777p 0.555588mV 618090.52p 0.556235mV 618107.358p 0.557275mV 618112.895p 0.557629mV 618124.492p 0.557984mV 619007.549p 0.548125mV 619011.843p 0.547736mV 619019.663p 0.546983mV 619031.311p 0.543264mV 621004.334p 0.547764mV 621004.635p 0.547764mV 621010.287p 0.547406mV 621042.647p 0.548517mV 621050.722p 0.549617mV 621053.447p 0.549617mV 621074.395p 0.551816mV 621082.747p 0.555115mV 621090.861p 0.559882mV 622021.236p 0.553422mV 622026.983p 0.553388mV 622073.052p 0.562189mV 623003.179p 0.554023mV 623039.721p 0.553062mV 623042.177p 0.552615mV 623043.85p 0.552615mV 623053.115p 0.550626mV 623067.591p 0.547098mV 623074.349p 0.545922mV 623077.577p 0.54511mV 623081.553p 0.544663mV 623114.845p 0.544509mV 623148.074p 0.547869mV 623155.066p 0.550237mV 623173.178p 0.55288mV 623177.895p 0.553521mV 623194.417p 0.556191mV 624033.14p 0.554013mV 624038.163p 0.553246mV 624070.959p 0.554461mV 624091.44p 0.557249mV 624109.42p 0.558991mV 624109.471p 0.558991mV 625014.185p 0.553373mV 625022.473p 0.553592mV 625027.609p 0.554249mV 625031.587p 0.555271mV 625039.911p 0.556658mV 625041.657p 0.55841mV 625047.421p 0.559798mV 626007.3p 0.546404mV 626050.565p 0.551086mV 626055.673p 0.552462mV 626065.773p 0.556318mV 627006.03p 0.554218mV 627021.905p 0.55509mV 627027.099p 0.555136mV 627028.758p 0.555136mV 627029.896p 0.555136mV 627038.004p 0.554861mV 627047.638p 0.555316mV 627083.795p 0.560753mV 627092.957p 0.56195mV 627104.182p 0.562426mV 627105.297p 0.562484mV 627122.63p 0.562678mV 627140.558p 0.561519mV 627160.937p 0.559684mV 627173.291p 0.559518mV 627187.063p 0.55656mV 627217.271p 0.550394mV 627233.091p 0.547187mV 628008.32p 0.553292mV 628040.158p 0.548606mV 628067.186p 0.543261mV 629025.617p 0.543483mV 630019.563p 0.554559mV 630024.448p 0.554896mV 630037.268p 0.558105mV 630043.492p 0.559907mV 631002.949p 0.552785mV 631012.557p 0.552286mV 631023.895p 0.551784mV 631041.558p 0.553698mV 631053.974p 0.556846mV 631054.411p 0.556846mV 631075.825p 0.566745mV 632022.976p 0.553025mV 632034.937p 0.554146mV 632056.709p 0.552007mV 632088.897p 0.548759mV 633007.015p 0.546557mV 633010.042p 0.546235mV 633016.106p 0.545547mV 633019.934p 0.545547mV 633035.318p 0.542064mV 633053.861p 0.53853mV 634064.88p 0.553302mV 634082.165p 0.552687mV 635011.697p 0.546968mV 635023.816p 0.546754mV 635030.448p 0.545079mV 635051.153p 0.539529mV 635069.535p 0.537904mV 635078.397p 0.536194mV 636067.88p 0.541499mV 637011.789p 0.54862mV 637030.351p 0.546371mV 637042.968p 0.543778mV 637068.336p 0.541456mV 637091.435p 0.542331mV 638014.337p 0.549208mV 638015.373p 0.54923mV 638031.646p 0.547105mV 638047.224p 0.543882mV 638066.977p 0.537371mV 638068.447p 0.537371mV 639020.166p 0.548901mV 639044.254p 0.551145mV 639063.039p 0.555599mV 640011.849p 0.550068mV 640046.253p 0.554301mV 640054.942p 0.555329mV 640059.881p 0.556725mV 640068.405p 0.56062mV 641004.741p 0.549058mV 641005.807p 0.54907mV 641067.983p 0.555127mV 641075.035p 0.553365mV 641092.497p 0.552019mV 641101.946p 0.552472mV 642004.777p 0.549903mV 642022.897p 0.549129mV 642044.27p 0.551271mV 642062.373p 0.55487mV 642080.228p 0.552633mV 642119.328p 0.546342mV 643009.896p 0.550064mV 643010.587p 0.550361mV 643041.394p 0.556194mV 644012.068p 0.552274mV 644039.643p 0.552263mV 644054.035p 0.550787mV 644099.814p 0.552154mV 644111.977p 0.553562mV 644161.273p 0.557357mV 644185.072p 0.555756mV 644203.014p 0.557114mV 644233.504p 0.560125mV 644234.052p 0.560125mV 644238.844p 0.560801mV 644243.478p 0.561839mV 644252.32p 0.563541mV 644281.057p 0.567845mV 645016.039p 0.548161mV 645051.931p 0.542463mV 646009.589p 0.546294mV 646021.847p 0.546181mV 646045.37p 0.541611mV 646067.686p 0.53487mV 647006.693p 0.552089mV 647032.855p 0.549551mV 647059.513p 0.551033mV 647061.158p 0.551402mV 647072.948p 0.552508mV 647086.639p 0.552161mV 647124.626p 0.556634mV 647133.219p 0.558506mV 647138.822p 0.559264mV 648007.244p 0.552259mV 648046.102p 0.543966mV 649021.388p 0.55126mV 649109.302p 0.552962mV 649130.272p 0.548819mV 649154.681p 0.544312mV 649155.001p 0.543545mV 649159.532p 0.543545mV 650009.041p 0.550859mV 650034.4p 0.549895mV 650038.24p 0.549187mV 650055.954p 0.550001mV 650063.551p 0.551114mV 650079.097p 0.554448mV 650081.298p 0.556289mV 650084.674p 0.556289mV 650085.556p 0.558496mV 651002.015p 0.550959mV 651022.012p 0.551072mV 652000.272p 0.553359mV 652001.175p 0.553359mV 652006.14p 0.553327mV 652018.095p 0.552896mV 654022.187p 0.550845mV 654033.005p 0.552829mV 654055.435p 0.559832mV 654058.427p 0.559832mV 655008.606p 0.55428mV 655018.998p 0.553883mV 655023.405p 0.554234mV 655043.543p 0.552719mV 655063.3p 0.553407mV 655065.977p 0.554129mV 655078.177p 0.555209mV 656030.886p 0.553919mV 657001.936p 0.552921mV 657006.207p 0.552944mV 657019.165p 0.551896mV 657050.067p 0.546954mV 657051.428p 0.546954mV 657067.773p 0.54592mV 657087.432p 0.54305mV 658011.636p 0.552368mV 658033.095p 0.550964mV 658074.616p 0.546671mV 658079.188p 0.545215mV 659026.856p 0.553455mV 659054.892p 0.557863mV 659077.362p 0.55758mV 659099.129p 0.553756mV 659107.518p 0.551128mV 659112.68p 0.549268mV 659121.862p 0.544456mV 659141.213p 0.531172mV 660042.741p 0.547492mV 660082.948p 0.548098mV 660111.713p 0.55566mV 661013.613p 0.549816mV 661016.648p 0.549755mV 661024.35p 0.550058mV 661054.736p 0.547839mV 661064.819p 0.548065mV 661080.935p 0.552889mV 661103.861p 0.559172mV 662015.732p 0.552985mV 662041.525p 0.553143mV 662041.603p 0.553143mV 662057.964p 0.551936mV 662071.543p 0.549641mV 662107.913p 0.541739mV 662138.1p 0.533083mV 662139.203p 0.533083mV 662139.514p 0.533083mV 663012.273p 0.546092mV 663049.969p 0.550546mV 663057.12p 0.553979mV 664001.724p 0.551689mV 664007.087p 0.55161mV 664042.059p 0.541511mV 665052.952p 0.555652mV 665067.001p 0.552208mV 665071.865p 0.551064mV 665072.12p 0.551064mV 665088.466p 0.546907mV 665103.869p 0.542388mV 665104.636p 0.542388mV 665121.027p 0.540738mV 665135.864p 0.538022mV 665168.762p 0.532169mV 666011.063p 0.550473mV 666016.434p 0.550403mV 666017.497p 0.550403mV 666055.186p 0.549821mV 666091.035p 0.542669mV 667017.669p 0.547242mV 668031.305p 0.549746mV 668131.996p 0.541949mV 668179.766p 0.545993mV 669016.381p 0.5533mV 669037.845p 0.554527mV 669045.122p 0.556968mV 670047.928p 0.540915mV 670071.035p 0.538661mV 670094.103p 0.540429mV 670105.404p 0.540431mV 671001.938p 0.548066mV 671013.408p 0.548282mV 671025.195p 0.548431mV 671034.033p 0.547994mV 671039.123p 0.547193mV 671124.944p 0.543658mV 672009.489p 0.547024mV 672014.877p 0.547416mV 672041.222p 0.553057mV 672042.77p 0.553057mV 672046.251p 0.555279mV 673012.432p 0.551721mV 673028.524p 0.550693mV 673029.855p 0.550693mV 673031.651p 0.550348mV 673033.668p 0.550348mV 673039.548p 0.549634mV 673042.377p 0.549285mV 673085.719p 0.546369mV 674010.419p 0.554657mV 674012.034p 0.554657mV 674039.161p 0.55191mV 674065.374p 0.542985mV 674070.506p 0.541187mV 675007.71p 0.550753mV 675022.88p 0.551582mV 675076.079p 0.561748mV 675094.842p 0.566228mV 676063.03p 0.546834mV 676071.09p 0.547287mV 676087.273p 0.550686mV 676094.034p 0.551813mV 676105.023p 0.553721mV 676128.418p 0.558188mV 676143.298p 0.560427mV 676148.318p 0.56044mV 676154.383p 0.560817mV 676157.159p 0.560827mV 676168.922p 0.560475mV 676169.181p 0.560475mV 676187.913p 0.560471mV 677030.4p 0.545962mV 677039.087p 0.54529mV 677052.719p 0.544726mV 677069.281p 0.54378mV 677084.98p 0.541716mV 677087.572p 0.541022mV 677090.618p 0.54069mV 678006.73p 0.552917mV 678007.265p 0.552917mV 678025.82p 0.553464mV 678030.764p 0.553784mV 678031.216p 0.553784mV 678053.397p 0.555071mV 678066.722p 0.55824mV 678087.084p 0.560302mV 678153.607p 0.554855mV 678162.282p 0.552379mV 679001.073p 0.552748mV 679056.228p 0.552053mV 679061.841p 0.551583mV 679066.054p 0.551478mV 679071.879p 0.551006mV 679089.107p 0.547383mV 679093.142p 0.54544mV 680001.354p 0.546498mV 680013.545p 0.546967mV 680071.25p 0.550576mV 680109.221p 0.550711mV 680133.825p 0.55078mV 680134.305p 0.55078mV 681037.502p 0.553735mV 682000.485p 0.550315mV 682016.766p 0.550446mV 682033.294p 0.550209mV 682034.316p 0.550209mV 682072.298p 0.548102mV 682073.176p 0.548102mV 682080.704p 0.54757mV 682084.616p 0.54757mV 682096.337p 0.547678mV 682099.123p 0.547678mV 682102.094p 0.547223mV 682104.173p 0.547223mV 682113.383p 0.545945mV 682130.069p 0.545559mV 682130.489p 0.545559mV 682145.27p 0.544146mV 682148.809p 0.544146mV 683005.797p 0.55033mV 683007.021p 0.55033mV 683029.002p 0.551736mV 683049.23p 0.556085mV 683052.087p 0.557908mV 684002.021p 0.545688mV 684026.041p 0.548265mV 684055.18p 0.552011mV 684064.923p 0.553186mV 684094.055p 0.561377mV 685009.155p 0.546443mV 685028.413p 0.546286mV 685031.609p 0.54588mV 685084.016p 0.549461mV 685098.062p 0.552617mV 685145.319p 0.554856mV 685147.53p 0.554856mV 685158.501p 0.553732mV 685201.868p 0.546804mV 685214.826p 0.54574mV 686038.963p 0.544895mV 686039.111p 0.544895mV 686049.731p 0.542466mV 686079.127p 0.538779mV 687023.471p 0.551549mV 687048.615p 0.550774mV 687064.527p 0.547084mV 687081.609p 0.544088mV 687082.768p 0.544088mV 687083.341p 0.544088mV 688022.228p 0.550093mV 688054.148p 0.545703mV 688059.908p 0.545028mV 688065.772p 0.543303mV 688078.283p 0.543027mV 689007.533p 0.550438mV 689027.819p 0.547727mV 689038.746p 0.545268mV 690017.347p 0.549698mV 690064.258p 0.544689mV 690068.493p 0.544655mV 690070.181p 0.544254mV 690079.784p 0.544218mV 690081.04p 0.543814mV 690090.719p 0.542636mV 690101.014p 0.542912mV 690106.301p 0.543595mV 690115.172p 0.54532mV 690126.516p 0.547769mV 690133.212p 0.54954mV 690186.115p 0.566156mV 691016.021p 0.554459mV 692020.227p 0.553747mV 692074.08p 0.560375mV 692080.96p 0.55854mV 692094.48p 0.557456mV 692104.019p 0.555663mV 694000.478p 0.547352mV 694008.872p 0.547433mV 694010.367p 0.547148mV 694016.988p 0.546495mV 694022.534p 0.546207mV 695002.548p 0.547364mV 695034.774p 0.546963mV 695074.161p 0.545374mV 695077.077p 0.544617mV 695083.918p 0.543492mV 696003.114p 0.552226mV 696022.358p 0.551784mV 696052.562p 0.549665mV 696055.203p 0.548275mV 697015.477p 0.546703mV 697023.314p 0.547055mV 697063.1p 0.55139mV 697081.699p 0.554352mV 698032.465p 0.543168mV 699009.258p 0.554671mV 699042.669p 0.545543mV 699042.901p 0.545543mV 700004.814p 0.554238mV 700028.56p 0.552882mV 700030.802p 0.551804mV 700032.568p 0.551804mV 701008.791p 0.547674mV 701012.379p 0.547949mV 701099.129p 0.548492mV 701105.339p 0.54865mV 701109.126p 0.54865mV 702010.207p 0.546611mV 702014.798p 0.546611mV 702016.098p 0.545921mV 702024.423p 0.544865mV 702056.291p 0.546967mV 702068.299p 0.548869mV 702071.461p 0.550004mV 703063.584p 0.55543mV 703078.013p 0.556616mV 703111.387p 0.558378mV 703123.601p 0.560321mV 704022.17p 0.547568mV 704034.953p 0.547198mV 704047.463p 0.543909mV 705045.557p 0.552061mV 705074.109p 0.552195mV 705076.072p 0.552299mV 705099.592p 0.549072mV 705123.206p 0.544138mV 705128.816p 0.544246mV 705243.278p 0.549168mV 705254.54p 0.551291mV 706008.591p 0.552503mV 706013.677p 0.552866mV 706078.487p 0.553648mV 706078.841p 0.553648mV 706126.369p 0.551298mV 706143.106p 0.552133mV 706164.558p 0.553773mV 707002.267p 0.545928mV 707026.81p 0.545503mV 707082.337p 0.552701mV 708000.666p 0.553735mV 708024.797p 0.55466mV 708053.604p 0.559685mV 708062.281p 0.560874mV 708070.97p 0.561335mV 708087.693p 0.560392mV 708091.32p 0.559348mV 708096.775p 0.558672mV 708107.792p 0.557686mV 708109.146p 0.557686mV 708163.907p 0.547239mV 709020.328p 0.552693mV 709022.771p 0.552693mV 709049.837p 0.548345mV 709053.313p 0.54725mV 709065.28p 0.544674mV 710002.431p 0.548124mV 710009.13p 0.548057mV 710017.792p 0.546831mV 710018.159p 0.546831mV 710041.111p 0.54396mV 710041.638p 0.54396mV 710042.875p 0.54396mV 710095.417p 0.541425mV 710110.58p 0.541215mV 710129.373p 0.540636mV 710131.135p 0.540198mV 710172.279p 0.546913mV 710180.152p 0.548597mV 711038.354p 0.551711mV 711055.97p 0.556288mV 711080.877p 0.567142mV 712007.487p 0.545809mV 712022.028p 0.547748mV 712032.637p 0.548681mV 712042.982p 0.54889mV 712043.94p 0.54889mV 712069.742p 0.548544mV 712118.201p 0.53525mV 712121.027p 0.533378mV 712207.672p 0.523718mV 712267.265p 0.524527mV 713038.989p 0.559904mV 713041.489p 0.561775mV 714016.151p 0.546572mV 714022.431p 0.546857mV 714037.745p 0.547709mV 714040.775p 0.547261mV 714050.672p 0.547465mV 714066.461p 0.548321mV 714096.33p 0.555544mV 714098.203p 0.555544mV 715040.139p 0.552157mV 715058.54p 0.547982mV 716004.802p 0.549948mV 716012.792p 0.550461mV 716036.654p 0.554493mV 716039.656p 0.554493mV 717004.851p 0.553313mV 717026.936p 0.553036mV 717031.975p 0.55203mV 717046.722p 0.547547mV 717047.991p 0.547547mV 718013.459p 0.545844mV 718023.715p 0.546284mV 718025.626p 0.547052mV 718060.936p 0.557556mV 719002.22p 0.549844mV 719002.388p 0.549844mV 719026.936p 0.5467mV 719031.77p 0.546287mV 719060.503p 0.547782mV 719061.862p 0.547782mV 720013.568p 0.55008mV 720024.898p 0.550324mV 720034.329p 0.549839mV 720079.035p 0.539799mV 721011.584p 0.545829mV 721018.98p 0.545763mV 721022.51p 0.546062mV 721023.888p 0.546062mV 721027.581p 0.545993mV 721039.939p 0.544756mV 722012.841p 0.548136mV 722043.399p 0.553684mV 722069.499p 0.558899mV 722071.152p 0.559296mV 723006.609p 0.551668mV 723031.02p 0.548405mV 723035.933p 0.547674mV 723037.792p 0.547674mV 723039.775p 0.547674mV 724001.007p 0.550884mV 724041.035p 0.546456mV 724043.985p 0.546456mV 724047.326p 0.544984mV 724060.649p 0.542746mV 724063.481p 0.542746mV 724072.219p 0.540872mV 725024.47p 0.552521mV 725025.953p 0.553258mV 725041.212p 0.555478mV 725062.216p 0.556275mV 725083.115p 0.554193mV 725096.524p 0.553939mV 726011.971p 0.548316mV 726033.111p 0.553381mV 726036.801p 0.554831mV 726059.286p 0.559922mV 727031.959p 0.553602mV 727044.596p 0.553068mV 727055.227p 0.551714mV 727061.602p 0.550529mV 727082.66p 0.542846mV 728025.347p 0.552803mV 728063.498p 0.550149mV 728065.832p 0.549353mV 728082.009p 0.546965mV 728109.82p 0.542973mV 728123.938p 0.542021mV 728137.202p 0.540683mV 728145.839p 0.541604mV 728164.431p 0.543513mV 728179.6p 0.545768mV 728189.557p 0.547384mV 728191.713p 0.548372mV 728219.518p 0.554398mV 728258.442p 0.568897mV 729013.704p 0.55207mV 729035.719p 0.554014mV 729041.313p 0.554331mV 729100.434p 0.542876mV 730012.028p 0.553533mV 730040.707p 0.548232mV 731030.142p 0.553287mV 731051.132p 0.551035mV 731080.339p 0.545446mV 731097.821p 0.541344mV 731098.664p 0.541344mV 732002.96p 0.552042mV 732010.248p 0.552533mV 732048.986p 0.558474mV 732055.306p 0.560447mV 733000.437p 0.551385mV 733016.322p 0.550951mV 733043.883p 0.548275mV 733051.616p 0.546397mV 733064.545p 0.543781mV 733079.654p 0.541851mV 733091.501p 0.539526mV 734000.422p 0.553614mV 734051.593p 0.550419mV 734089.538p 0.549237mV 734094.805p 0.548846mV 735030.409p 0.547861mV 735057.314p 0.551534mV 736012.355p 0.552009mV 736025.328p 0.554629mV 736030.406p 0.555749mV 736034.453p 0.555749mV 736036.685p 0.557238mV 737033.516p 0.545907mV 737034.316p 0.545907mV 737057.848p 0.539965mV 737073.815p 0.536974mV 737078.771p 0.535485mV 737085.347p 0.532132mV 738001.091p 0.547095mV 738004.01p 0.547095mV 738016.288p 0.546265mV 738071.867p 0.545633mV 738071.889p 0.545633mV 738088.039p 0.544703mV 738093.347p 0.544387mV 738094.226p 0.544387mV 738099.121p 0.544432mV 738101.532p 0.544107mV 739009.49p 0.547481mV 739010.809p 0.547066mV 739045.591p 0.547065mV 739067.538p 0.54537mV 739073.446p 0.544943mV 739096.477p 0.546068mV 739106.838p 0.547746mV 739107.127p 0.547746mV 739108.508p 0.547746mV 739156.951p 0.561176mV 739168.883p 0.563572mV 739173.656p 0.56459mV 739181.552p 0.567mV 739184.98p 0.567mV 740027.795p 0.552977mV 740053.149p 0.550789mV 741049.501p 0.557761mV 741054.882p 0.558966mV 742000.974p 0.546768mV 742003.144p 0.546768mV 743010.14p 0.552297mV 743057.668p 0.552367mV 743061.96p 0.551205mV 743084.93p 0.549495mV 743092.462p 0.549013mV 743092.6p 0.549013mV 743143.539p 0.54227mV 743150.816p 0.540342mV 743160.251p 0.536953mV 743166.996p 0.534709mV 743196.709p 0.523045mV 743198.569p 0.523045mV 744001.696p 0.548782mV 744011.399p 0.549168mV 744032.014p 0.551405mV 744047.99p 0.553271mV 744053.6p 0.553652mV 744060.376p 0.555517mV 745006.778p 0.553831mV 745013.85p 0.553507mV 745050.175p 0.553776mV 745056.975p 0.555262mV 745058.394p 0.555262mV 745085.102p 0.564523mV 745086.084p 0.564523mV 745103.714p 0.567515mV 745104.716p 0.567515mV 745112.675p 0.568667mV 745131.149p 0.573196mV 746007.5p 0.553926mV 746018.044p 0.553712mV 746057.369p 0.557954mV 746064.922p 0.558392mV 746081.811p 0.560881mV 746142.663p 0.567053mV 746153.135p 0.569096mV 747007.851p 0.55352mV 747011.111p 0.553158mV 747080.242p 0.559483mV 747095.553p 0.56065mV 747107.844p 0.561083mV 747108.969p 0.561083mV 748000.231p 0.551929mV 748007.035p 0.552014mV 748013.882p 0.551734mV 748015.592p 0.551819mV 748030.203p 0.553541mV 748047.459p 0.554902mV 748085.364p 0.563003mV 749022.972p 0.549057mV 749029.232p 0.550582mV 749047.136p 0.557437mV 750070.748p 0.554659mV 750083.278p 0.553754mV 750129.208p 0.551682mV 750129.999p 0.551682mV 750134.267p 0.551408mV 750140.37p 0.551223mV 750143.655p 0.551223mV 750166.489p 0.55019mV 750182.55p 0.547503mV 750187.858p 0.546846mV 750196.073p 0.545158mV 751001.3p 0.551099mV 751019.349p 0.550006mV 751028.403p 0.54964mV 751042.041p 0.548169mV 751042.56p 0.548169mV 751069.308p 0.547392mV 752003.663p 0.547094mV 753006.384p 0.546028mV 753036.685p 0.544217mV 753064.342p 0.548236mV 753085.71p 0.553355mV 754001.287p 0.553107mV 754012.645p 0.552582mV 754018.388p 0.552502mV 754042.203p 0.554645mV 754062.449p 0.555768mV 754075.829p 0.557347mV 754100.504p 0.557321mV 754101.567p 0.557321mV 754111.052p 0.557541mV 754112.995p 0.557541mV 754141.504p 0.557522mV 755022.818p 0.554578mV 755038.71p 0.557073mV 756007.154p 0.553102mV 756038.594p 0.557294mV 756043.154p 0.559152mV 756043.187p 0.559152mV 756059.954p 0.564001mV 757000.53p 0.551493mV 757013.779p 0.551908mV 757017.496p 0.552665mV 757041.924p 0.558297mV 757047.04p 0.559065mV 758018.299p 0.549909mV 758051.085p 0.557561mV 759002.956p 0.549844mV 759021.494p 0.549573mV 759022.978p 0.549573mV 759032.019p 0.548345mV 759032.057p 0.548345mV 759048.813p 0.547789mV 759060.219p 0.545408mV 759071.475p 0.541992mV 759074.324p 0.541992mV 759076.717p 0.539735mV 759084.058p 0.537842mV 760009.855p 0.548966mV 760012.329p 0.549272mV 760039.386p 0.55046mV 760066.143p 0.550564mV 760071.61p 0.550165mV 760089.903p 0.548255mV 760136.418p 0.533867mV 760136.762p 0.533867mV 760148.791p 0.529827mV 761005.344p 0.553646mV 761043.708p 0.555205mV 761059.975p 0.560428mV 762019.125p 0.549418mV 762049.99p 0.554663mV 762069.74p 0.561594mV 763013.299p 0.551693mV 763026.84p 0.551076mV 763033.517p 0.551358mV 763043.392p 0.553021mV 763068.322p 0.554819mV 763076.717p 0.55577mV 763094.543p 0.557032mV 763121.523p 0.551244mV 763121.578p 0.551244mV 763145.291p 0.540832mV 763155.443p 0.536745mV 763172.78p 0.530791mV 763183.72p 0.526689mV 763184.365p 0.526689mV 763192.192p 0.523305mV 764035.445p 0.547896mV 764041.821p 0.54602mV 764046.991p 0.543777mV 764067.369p 0.538443mV 764075.548p 0.537946mV 766026.02p 0.546264mV 766067.476p 0.538942mV 767013.786p 0.551616mV 767016.287p 0.551565mV 767038.853p 0.550622mV 767055.491p 0.548935mV 767082.162p 0.546053mV 767083.762p 0.546053mV 768032.724p 0.554374mV 768073.719p 0.552473mV 768116.303p 0.552806mV 768135.095p 0.551957mV 768158.102p 0.545306mV 768171.222p 0.538693mV 768175.499p 0.535758mV 768185.329p 0.529522mV 768204.424p 0.522163mV 769001.393p 0.549933mV 769020.033p 0.548257mV 769023.541p 0.548257mV 769088.53p 0.546846mV 769094.053p 0.547158mV 769099.212p 0.547836mV 769100.946p 0.548149mV 769106.561p 0.548829mV 769136.402p 0.556966mV 770003.309p 0.550142mV 770033.287p 0.550127mV 771005.307p 0.55453mV 771012.967p 0.554179mV 771037.619p 0.548388mV 771038.757p 0.548388mV 771049.698p 0.545838mV 772004.148p 0.554396mV 772017.161p 0.555221mV 772033.019p 0.557139mV 772050.926p 0.55897mV 772086.834p 0.560964mV 772089.031p 0.560964mV 773014.82p 0.54665mV 773022.966p 0.547163mV 773026.124p 0.547967mV 773061.409p 0.552148mV 773085.276p 0.551098mV 773104.676p 0.553557mV 773117.715p 0.554936mV 773120.483p 0.555402mV 773124.091p 0.555402mV 774022.505p 0.547686mV 774060.721p 0.546929mV 774072.004p 0.549283mV 774079.645p 0.550642mV 774092.397p 0.556913mV 775005.784p 0.54885mV 775071.856p 0.544494mV 775090.951p 0.538303mV 775119.285p 0.537078mV 775133.446p 0.536734mV 776057.196p 0.552887mV 776088.134p 0.550671mV 776094.646p 0.549503mV 777013.217p 0.54788mV 777016.506p 0.547132mV 777100.512p 0.555071mV 777114.997p 0.559757mV 778018.886p 0.545877mV 778054.031p 0.54542mV 778069.8p 0.544428mV 778094.408p 0.542011mV 779019.831p 0.553544mV 779022.408p 0.553195mV 779024.038p 0.553195mV 780012.015p 0.549194mV 780023.497p 0.549695mV 780025.727p 0.550494mV 780036.873p 0.551728mV 780039.061p 0.551728mV 780042.676p 0.552162mV 780062.762p 0.556107mV 780063.758p 0.556107mV 780076.009p 0.557441mV 780090.643p 0.557705mV 781003.651p 0.546428mV 781019.461p 0.545151mV 781043.843p 0.53933mV 781054.129p 0.537346mV 782013.194p 0.546519mV 782042.686p 0.548216mV 782044.477p 0.548216mV 782079.443p 0.554342mV 783007.121p 0.552441mV 783008.043p 0.552441mV 783045.444p 0.553186mV 783089.262p 0.56488mV 784032.313p 0.55286mV 784052.012p 0.555117mV 786019.146p 0.552354mV 786037.676p 0.554124mV 786038.023p 0.554124mV 787006.941p 0.550643mV 787007.052p 0.550643mV 787014.196p 0.55034mV 787020.035p 0.548637mV 787024.435p 0.548637mV 787054.96p 0.545695mV 787074.955p 0.542956mV 788028.785p 0.547845mV 788029.831p 0.547845mV 788076.482p 0.53998mV 789009.296p 0.553088mV 789033.953p 0.553289mV 789063.55p 0.557814mV 789070.289p 0.560296mV 789098.807p 0.563056mV 789103.602p 0.562665mV 789105.359p 0.561911mV 789144.843p 0.558895mV 789149.093p 0.558159mV 789189.813p 0.545012mV 789202.751p 0.537701mV 789204.562p 0.537701mV 790060.466p 0.552503mV 790064.161p 0.552503mV 791006.228p 0.550507mV 791059.784p 0.550509mV 791078.852p 0.556509mV 791079.215p 0.556509mV 792035.351p 0.552107mV 792037.365p 0.552107mV 792040.555p 0.55183mV 792078.748p 0.555749mV 792085.506p 0.557028mV 792096.152p 0.559043mV 792113.41p 0.560801mV 793012.285p 0.547408mV 793043.456p 0.552024mV 794007.513p 0.545704mV 794010.167p 0.545984mV 794021.775p 0.546176mV 794080.32p 0.534121mV 796064.143p 0.553125mV 796123.612p 0.562196mV 796130.402p 0.563346mV 796143.943p 0.565232mV 796177.258p 0.564384mV 796220.369p 0.563678mV 796237.571p 0.564909mV 796246.594p 0.565365mV 796250.432p 0.565046mV 796251.871p 0.565046mV 796253.579p 0.565046mV 796257.475p 0.565093mV 796268.549p 0.564822mV 796310.653p 0.561998mV 796311.211p 0.561998mV 796350.45p 0.551436mV 797032.739p 0.54477mV 797039.067p 0.543966mV 797104.948p 0.548468mV 797148.403p 0.550807mV 797158.485p 0.549608mV 797172.366p 0.546553mV 797172.398p 0.546553mV 797174.381p 0.546553mV 797192.537p 0.53837mV 797223.947p 0.521707mV 798000.904p 0.552118mV 798012.853p 0.552423mV 798013.666p 0.552423mV 799008.855p 0.550989mV 799018.381p 0.550626mV 799021.425p 0.550261mV 799077.038p 0.554259mV 799080.721p 0.555353mV 799100.661p 0.558279mV 799125.762p 0.563457mV 800004.618p 0.5474mV 800047.269p 0.546317mV 800050.177p 0.546633mV 800052.038p 0.546633mV 800087.861p 0.553913mV 800110.194p 0.560552mV 800112.914p 0.560552mV 800133.252p 0.564714mV 800147.135p 0.570056mV 801007.111p 0.547237mV 801009.994p 0.547237mV 801029.891p 0.54599mV 802064.379p 0.553663mV 802075.569p 0.555811mV 802082.163p 0.556288mV 802084.98p 0.556288mV 802093.762p 0.55835mV 803015.208p 0.545645mV 803027.321p 0.546621mV 803033.591p 0.547656mV 804000.471p 0.551317mV 804008.899p 0.551265mV 804034.99p 0.547716mV 804052.0p 0.543111mV 805007.0p 0.551209mV 805026.565p 0.54764mV 805027.583p 0.54764mV 805031.431p 0.546564mV 806003.219p 0.548924mV 806005.015p 0.548868mV 806049.436p 0.546986mV 806052.163p 0.545838mV 806056.378p 0.545057mV 806060.2p 0.54391mV 806067.308p 0.542397mV 806075.103p 0.539002mV 807002.355p 0.550016mV 807025.246p 0.546301mV 807035.329p 0.543718mV 807040.01p 0.541875mV 807049.623p 0.540397mV 807056.764p 0.538528mV 807061.103p 0.538136mV 808016.374p 0.549398mV 808021.866p 0.549768mV 808088.765p 0.549826mV 808093.527p 0.549466mV 808132.896p 0.536321mV 809021.559p 0.553807mV 809039.25p 0.552987mV 809062.165p 0.553832mV 809088.761p 0.5558mV 809090.158p 0.555541mV 809092.471p 0.555541mV 809113.77p 0.555992mV 809125.412p 0.55307mV 809135.498p 0.551502mV 809148.699p 0.550674mV 809213.388p 0.546453mV 810030.493p 0.548177mV 810041.225p 0.547824mV 810045.597p 0.547831mV 810057.953p 0.546747mV 810079.078p 0.543111mV 810085.346p 0.541286mV 811007.511p 0.552387mV 811015.809p 0.553584mV 811061.245p 0.551553mV 811064.803p 0.551553mV 811076.842p 0.546268mV 811081.029p 0.543775mV 812001.956p 0.55392mV 812005.197p 0.553959mV 812012.234p 0.554365mV 812023.047p 0.55408mV 812035.79p 0.554574mV 812039.829p 0.554574mV 812061.096p 0.552978mV 812074.55p 0.551247mV 812114.95p 0.547983mV 812117.133p 0.5473mV 812132.288p 0.544513mV 813010.616p 0.546605mV 813104.481p 0.540432mV 813110.549p 0.54065mV 813111.534p 0.54065mV 813129.614p 0.543717mV 814007.763p 0.548078mV 814022.083p 0.548797mV 814030.288p 0.550621mV 814041.643p 0.55245mV 814050.12p 0.553556mV 814058.443p 0.554296mV 815008.45p 0.54649mV 815010.659p 0.546902mV 815056.003p 0.552493mV 815072.225p 0.552694mV 815122.94p 0.548847mV 815144.811p 0.547122mV 816025.159p 0.550014mV 816067.118p 0.551823mV 817006.617p 0.552031mV 817023.981p 0.554349mV 817059.048p 0.552885mV 817059.96p 0.552885mV 817064.774p 0.55185mV 817071.598p 0.550882mV 817111.96p 0.543399mV 817113.528p 0.543399mV 817229.789p 0.535489mV 817230.355p 0.535151mV 817263.349p 0.534885mV 818026.55p 0.551303mV 818040.661p 0.557662mV 819005.695p 0.550152mV 819036.226p 0.555856mV 819066.283p 0.555042mV 819071.192p 0.555464mV 819091.864p 0.558641mV 819093.8p 0.558641mV 819095.96p 0.559444mV 820002.237p 0.549849mV 820027.209p 0.550239mV 820033.791p 0.55127mV 820041.367p 0.552969mV 820056.425p 0.55608mV 820082.531p 0.556215mV 821018.484p 0.550861mV 821029.955p 0.552041mV 821049.738p 0.55733mV 822000.615p 0.546463mV 822018.18p 0.545469mV 822032.31p 0.541913mV 822040.232p 0.540145mV 823009.256p 0.551336mV 823052.597p 0.543664mV 824000.397p 0.549554mV 824031.249p 0.549056mV 824056.67p 0.548176mV 825015.807p 0.552021mV 825033.307p 0.553617mV 825043.426p 0.554806mV 825060.563p 0.553542mV 825095.326p 0.554309mV 825127.612p 0.55216mV 825138.874p 0.549752mV 825150.204p 0.545601mV 825150.691p 0.545601mV 825179.035p 0.535757mV 825201.044p 0.530603mV 825217.466p 0.529651mV 826039.808p 0.552424mV 826042.048p 0.55274mV 826047.786p 0.552689mV 826070.152p 0.556451mV 826070.915p 0.556451mV 826096.617p 0.563516mV 827013.991p 0.553557mV 827028.613p 0.553973mV 827045.386p 0.556964mV 827072.831p 0.560353mV 827094.708p 0.560468mV 828035.129p 0.550437mV 828040.461p 0.549979mV 828049.197p 0.549156mV 828050.078p 0.547966mV 828050.94p 0.547966mV 828069.285p 0.546584mV 828094.327p 0.549371mV 828095.897p 0.549998mV 828149.272p 0.544174mV 828162.393p 0.543824mV 828194.45p 0.542674mV 829038.226p 0.555371mV 829050.309p 0.554799mV 829093.572p 0.55448mV 830024.461p 0.550891mV 830043.078p 0.551993mV 830060.332p 0.552382mV 830069.583p 0.552483mV 830087.496p 0.553634mV 832000.756p 0.55095mV 832010.94p 0.551336mV 832063.198p 0.546727mV 832104.145p 0.54389mV 832111.772p 0.542798mV 832125.15p 0.539499mV 832138.222p 0.536918mV 833008.723p 0.553109mV 833033.506p 0.549893mV 833034.197p 0.549893mV 833041.104p 0.546619mV 834016.353p 0.553119mV 834040.611p 0.553083mV 834042.226p 0.553083mV 834074.898p 0.558116mV 834089.417p 0.561939mV 835000.69p 0.548423mV 835012.883p 0.54824mV 835026.201p 0.545949mV 835029.683p 0.545949mV 835047.757p 0.546288mV 835057.753p 0.545348mV 835088.13p 0.541734mV 836015.357p 0.553965mV 836023.614p 0.554403mV 836055.094p 0.559653mV 836078.125p 0.566535mV 837001.023p 0.551661mV 837003.211p 0.551661mV 837040.213p 0.551891mV 837067.224p 0.556712mV 837077.771p 0.559895mV 838005.921p 0.548994mV 838012.899p 0.548664mV 838037.857p 0.547376mV 838042.633p 0.547775mV 838051.693p 0.548938mV 838094.477p 0.554319mV 839028.243p 0.55107mV 839035.527p 0.555017mV 840029.384p 0.544765mV 840033.191p 0.545069mV 840037.796p 0.545738mV 840068.81p 0.551574mV 841017.846p 0.553338mV 841033.235p 0.549713mV 842023.339p 0.553677mV 842050.52p 0.559923mV 842054.205p 0.559923mV 843004.256p 0.554087mV 843017.405p 0.553129mV 843050.735p 0.549022mV 843051.136p 0.549022mV 843056.462p 0.549053mV 843063.088p 0.548715mV 843098.66p 0.550623mV 843112.14p 0.552782mV 844004.942p 0.552792mV 844005.23p 0.552845mV 844022.888p 0.551543mV 844023.821p 0.551543mV 844084.966p 0.544788mV 845002.188p 0.55296mV 845020.156p 0.553117mV 845055.81p 0.549311mV 845104.681p 0.553374mV 846053.123p 0.557738mV 846053.84p 0.557738mV 846081.966p 0.559263mV 846107.608p 0.559091mV 846147.284p 0.55024mV 846151.253p 0.549148mV 846153.671p 0.549148mV 846163.21p 0.547337mV 846166.691p 0.545888mV 846182.717p 0.540093mV 846185.93p 0.537921mV 846205.334p 0.530711mV 846215.509p 0.526012mV 846255.422p 0.50571mV 847026.983p 0.550364mV 847043.242p 0.546037mV 847047.507p 0.544593mV 847057.702p 0.542794mV 848005.437p 0.554357mV 848063.988p 0.563696mV 848065.017p 0.565223mV 849071.57p 0.539404mV 849072.743p 0.539404mV 849076.903p 0.538626mV 850003.968p 0.546478mV 850006.543p 0.54653mV 850037.3p 0.542087mV 851009.465p 0.553487mV 851021.676p 0.553324mV 851065.511p 0.557901mV 851097.381p 0.558636mV 851176.392p 0.565142mV 852017.034p 0.549623mV 852017.381p 0.549623mV 852033.157p 0.550291mV 852042.084p 0.549884mV 852046.093p 0.549131mV 852062.524p 0.54614mV 852091.894p 0.54414mV 852096.657p 0.544103mV 852106.832p 0.545117mV 852109.722p 0.545117mV 852137.771p 0.550286mV 852146.149p 0.554185mV 852154.837p 0.55595mV 852162.468p 0.559843mV 852169.238p 0.561242mV 852176.268p 0.564408mV 852205.177p 0.572496mV 852214.501p 0.573551mV 852216.634p 0.574975mV 853030.219p 0.55487mV 853050.187p 0.562191mV 853052.314p 0.562191mV 853055.248p 0.563662mV 854027.184p 0.543779mV 854035.016p 0.541091mV 854044.418p 0.539194mV 855002.713p 0.554183mV 855032.934p 0.553413mV 855037.615p 0.552732mV 855043.672p 0.552415mV 855045.244p 0.551732mV 855057.646p 0.551455mV 855063.883p 0.551861mV 855111.233p 0.551753mV 855123.865p 0.551398mV 856020.936p 0.550228mV 856023.388p 0.550228mV 856040.259p 0.548984mV 856072.106p 0.549672mV 856082.67p 0.548681mV 856119.13p 0.542074mV 856188.864p 0.552128mV 856190.198p 0.55321mV 856228.027p 0.559244mV 856243.191p 0.563503mV 856251.371p 0.567421mV 856281.63p 0.580564mV 856284.435p 0.580564mV 856306.988p 0.595545mV 856308.413p 0.595545mV 856325.732p 0.609141mV 856333.391p 0.612363mV 857012.179p 0.548295mV 857021.548p 0.547305mV 857045.925p 0.540258mV 858013.794p 0.547938mV 858038.161p 0.547547mV 858079.678p 0.543668mV 858088.037p 0.543415mV 859024.091p 0.548193mV 859067.934p 0.545577mV 859127.014p 0.531083mV 860005.32p 0.554454mV 860027.544p 0.552743mV 860046.006p 0.553228mV 860063.15p 0.555971mV 860087.618p 0.562278mV 861010.061p 0.552612mV 861036.401p 0.553789mV 861039.252p 0.553789mV 861047.903p 0.555066mV 861062.756p 0.558267mV 861089.252p 0.56315mV 861103.868p 0.564222mV 863005.859p 0.54526mV 863034.591p 0.54668mV 863035.241p 0.547329mV 864002.472p 0.553153mV 864032.343p 0.55874mV 864043.575p 0.56281mV 865001.403p 0.549336mV 865008.15p 0.549364mV 865016.953p 0.549052mV 865035.746p 0.550612mV 865065.899p 0.551836mV 865089.244p 0.554835mV 865096.169p 0.555238mV 865096.435p 0.555238mV 865098.578p 0.555238mV 865149.649p 0.563905mV 865151.733p 0.564311mV 865162.248p 0.566229mV 866034.13p 0.554373mV 866036.59p 0.555172mV 866036.809p 0.555172mV 866050.294p 0.559762mV 866069.716p 0.566185mV 866077.839p 0.570356mV 867007.665p 0.554624mV 867013.878p 0.554951mV 867035.883p 0.552556mV 867048.634p 0.550643mV 867049.008p 0.550643mV 867058.539p 0.550186mV 867067.441p 0.551185mV 867098.02p 0.552674mV 867100.442p 0.552246mV 867218.449p 0.561597mV 867221.289p 0.560388mV 868006.573p 0.552107mV 868012.961p 0.552479mV 868017.023p 0.552484mV 868031.61p 0.551774mV 868036.871p 0.551051mV 868048.526p 0.549239mV 868050.602p 0.54815mV 869026.509p 0.545864mV 869045.588p 0.544418mV 869046.607p 0.544418mV 869048.91p 0.544418mV 869053.206p 0.544053mV 869059.104p 0.543321mV 869079.979p 0.544026mV 869091.382p 0.548367mV 869095.908p 0.54981mV 869102.655p 0.551617mV 869115.506p 0.556306mV 869115.738p 0.556306mV 870010.953p 0.548777mV 870013.256p 0.548777mV 870084.463p 0.552401mV 870100.46p 0.549899mV 870106.646p 0.54909mV 870123.664p 0.547395mV 870147.125p 0.546254mV 870168.7p 0.545899mV 870176.464p 0.545346mV 870184.242p 0.544883mV 870186.738p 0.544053mV 871001.391p 0.550165mV 871011.778p 0.549831mV 871015.83p 0.549118mV 871019.275p 0.549118mV 871041.386p 0.54739mV 871044.783p 0.54739mV 871049.595p 0.547412mV 871056.881p 0.547823mV 871070.188p 0.545699mV 871086.486p 0.541015mV 871113.228p 0.53342mV 872024.69p 0.551209mV 872037.802p 0.547804mV 872055.862p 0.545445mV 872070.375p 0.546029mV 872103.867p 0.546769mV 872121.098p 0.547945mV 872154.664p 0.54999mV 872217.334p 0.577839mV 873001.57p 0.546465mV 873001.841p 0.546465mV 873027.874p 0.547858mV 873049.419p 0.547078mV 873053.598p 0.546701mV 873073.802p 0.543733mV 873089.107p 0.541137mV 873090.27p 0.540757mV 873095.453p 0.54001mV 873132.782p 0.53617mV 873138.799p 0.53613mV 874061.699p 0.554244mV 874111.955p 0.553669mV 874117.546p 0.553665mV 876019.036p 0.546428mV 876020.699p 0.546712mV 876032.496p 0.548379mV 877041.486p 0.552334mV 877045.56p 0.553134mV 877056.455p 0.555829mV 877070.219p 0.558227mV 877096.523p 0.560783mV 877099.378p 0.560783mV 877128.446p 0.564572mV 877164.188p 0.56677mV 878008.753p 0.546337mV 878014.503p 0.546048mV 878018.092p 0.545393mV 878062.219p 0.546471mV 878062.268p 0.546471mV 878088.927p 0.548355mV 878105.672p 0.547257mV 878140.632p 0.541367mV 878157.169p 0.542768mV 878188.899p 0.543766mV 879005.189p 0.55216mV 879013.285p 0.551811mV 879015.907p 0.551097mV 879050.233p 0.545394mV 879076.495p 0.538172mV 880022.409p 0.54773mV 880041.698p 0.543398mV 880052.718p 0.540854mV 881003.048p 0.550235mV 881007.756p 0.550215mV 881021.779p 0.55162mV 881022.882p 0.55162mV 881060.675p 0.552244mV 881075.96p 0.551867mV 881104.643p 0.553713mV 881105.482p 0.555186mV 882006.838p 0.552274mV 882014.646p 0.552572mV 882018.317p 0.552505mV 882066.827p 0.547137mV 882102.334p 0.537939mV 882108.872p 0.53641mV 883037.674p 0.552877mV 883051.124p 0.553002mV 883059.74p 0.553042mV 883063.73p 0.552715mV 883064.685p 0.552715mV 883073.708p 0.553155mV 883084.219p 0.55359mV 883110.306p 0.552666mV 883127.853p 0.550896mV 883137.259p 0.550553mV 884035.44p 0.551664mV 884096.527p 0.555496mV 884131.535p 0.561244mV 885011.878p 0.550887mV 885016.671p 0.550215mV 885025.819p 0.549236mV 885041.285p 0.547215mV 885072.011p 0.545692mV 886001.136p 0.552572mV 886011.234p 0.552114mV 886061.744p 0.546188mV 886064.408p 0.546188mV 886068.018p 0.546141mV 886081.958p 0.548187mV 886083.247p 0.548187mV 886097.16p 0.549858mV 886097.186p 0.549858mV 886116.985p 0.5555mV 886127.958p 0.558695mV 886131.474p 0.560479mV 887019.718p 0.552986mV 887031.712p 0.550965mV 887052.277p 0.546804mV 887056.509p 0.545395mV 887057.195p 0.545395mV 888005.708p 0.552849mV 889029.856p 0.547708mV 889054.235p 0.544023mV 889071.602p 0.545133mV 889114.636p 0.547963mV 889130.828p 0.550417mV 889144.731p 0.549804mV 889146.89p 0.549676mV 889161.149p 0.549275mV 889204.182p 0.558238mV 889208.741p 0.559519mV 889227.907p 0.565332mV 890003.414p 0.55274mV 890018.304p 0.551904mV 890043.6p 0.550487mV 890095.33p 0.55083mV 890101.751p 0.551241mV 890133.306p 0.560562mV 890134.87p 0.560562mV 890135.734p 0.562774mV 890151.411p 0.569396mV 890165.23p 0.577836mV 890185.421p 0.58959mV 891026.398p 0.554066mV 891030.443p 0.554485mV 891035.737p 0.554536mV 891061.672p 0.556609mV 891109.523p 0.561403mV 891113.518p 0.562544mV 891159.902p 0.57325mV 891169.152p 0.573757mV 891177.962p 0.572826mV 891182.703p 0.57255mV 891188.067p 0.571914mV 891224.628p 0.567606mV 892014.814p 0.545806mV 892070.034p 0.545698mV 892070.221p 0.545698mV 892079.343p 0.545021mV 893002.358p 0.554306mV 893016.673p 0.554483mV 893043.434p 0.555261mV 893045.22p 0.554466mV 893053.346p 0.554037mV 893062.389p 0.552081mV 893098.595p 0.549044mV 893124.06p 0.549012mV 893147.708p 0.54563mV 894004.31p 0.554468mV 894017.836p 0.555747mV 894023.738p 0.556174mV 894036.924p 0.556729mV 894041.107p 0.556429mV 894050.196p 0.554734mV 894073.901p 0.548426mV 895003.194p 0.548547mV 895040.613p 0.556892mV 895049.874p 0.559038mV 897008.531p 0.552351mV 897010.376p 0.552637mV 897027.129p 0.554966mV 897055.147p 0.559315mV 898004.029p 0.548437mV 898005.803p 0.548459mV 898010.124p 0.548114mV 898024.838p 0.548522mV 898044.996p 0.548602mV 898078.362p 0.552034mV 898102.168p 0.559111mV 898102.19p 0.559111mV 899057.977p 0.556396mV 899080.786p 0.56374mV 900019.652p 0.551741mV 900020.777p 0.5521mV 900031.442p 0.551724mV 900038.26p 0.551721mV 900055.049p 0.555381mV 902000.607p 0.546327mV 903020.711p 0.550647mV 903092.426p 0.544826mV 903096.917p 0.544102mV 904002.442p 0.554383mV 904012.505p 0.554577mV 904096.606p 0.54281mV 904098.869p 0.54281mV 905029.416p 0.54903mV 905067.284p 0.545544mV 905077.342p 0.544306mV 905093.774p 0.543356mV 905142.022p 0.542885mV 906003.372p 0.548652mV 906012.196p 0.548345mV 906019.109p 0.548373mV 906164.011p 0.557963mV 907022.317p 0.552766mV 907046.038p 0.552431mV 907049.496p 0.552431mV 907050.702p 0.551995mV 907055.524p 0.551924mV 907084.443p 0.550453mV 907108.083p 0.550028mV 907113.67p 0.551031mV 907149.087p 0.559443mV 908012.593p 0.548048mV 908023.58p 0.549212mV 908031.917p 0.550376mV 908076.437p 0.546322mV 908105.664p 0.543237mV 908106.014p 0.543237mV 908132.129p 0.540793mV 908145.141p 0.539728mV 908154.216p 0.538635mV 909026.108p 0.545708mV 909034.808p 0.545268mV 909047.922p 0.545409mV 909115.815p 0.555703mV 909122.873p 0.556738mV 909124.342p 0.556738mV 910015.464p 0.548088mV 910023.621p 0.547778mV 910036.745p 0.548303mV 910061.826p 0.545978mV 910062.123p 0.545978mV 910067.149p 0.545287mV 910077.416p 0.543532mV 911022.877p 0.552586mV 911029.468p 0.553373mV 911033.157p 0.554527mV 911040.018p 0.556468mV 911081.741p 0.561375mV 911103.277p 0.556596mV 911135.574p 0.545944mV 911155.463p 0.543416mV 911204.075p 0.532891mV 911225.018p 0.531036mV 911276.876p 0.533947mV 911321.151p 0.545216mV 911331.758p 0.547723mV 911362.36p 0.555901mV 911369.861p 0.557315mV 911370.233p 0.559091mV 911372.062p 0.559091mV 911441.291p 0.585518mV 911468.479p 0.597492mV 911479.162p 0.60424mV 911520.782p 0.625614mV 911530.532p 0.626504mV 911540.593p 0.625927mV 912004.436p 0.546084mV 912004.992p 0.546084mV 912023.702p 0.545099mV 912027.446p 0.544305mV 912030.261p 0.543877mV 912058.103p 0.546489mV 912060.406p 0.547524mV 912065.286p 0.548926mV 912091.474p 0.551947mV 913011.186p 0.554417mV 914016.487p 0.550528mV 914022.46p 0.549482mV 914030.951p 0.547752mV 914057.426p 0.547948mV 914090.881p 0.558322mV 915002.32p 0.549663mV 915029.339p 0.54764mV 915050.994p 0.540116mV 915053.155p 0.540116mV 916008.789p 0.550975mV 916020.12p 0.5526mV 916067.563p 0.56116mV 916068.426p 0.56116mV 916068.963p 0.56116mV 917000.664p 0.547575mV 917058.574p 0.550272mV 917059.03p 0.550272mV 917076.144p 0.554973mV 917081.672p 0.55542mV 917084.973p 0.55542mV 917101.984p 0.558698mV 917122.226p 0.557649mV 918001.808p 0.55015mV 918023.103p 0.547659mV 918058.61p 0.538703mV 918067.79p 0.535967mV 919015.824p 0.551388mV 919023.561p 0.552458mV 919027.075p 0.553163mV 919041.595p 0.555293mV 919049.766p 0.556009mV 920002.497p 0.550034mV 920032.28p 0.555345mV 920042.273p 0.558104mV 921011.499p 0.552612mV 921026.418p 0.555863mV 921039.399p 0.559128mV 922007.965p 0.55164mV 923000.374p 0.549253mV 923030.768p 0.552244mV 923055.611p 0.561512mV 925001.123p 0.547701mV 925004.494p 0.547701mV 925061.167p 0.550079mV 925068.308p 0.550098mV 925100.673p 0.549518mV 925104.395p 0.549518mV 925107.228p 0.549542mV 925107.923p 0.549542mV 925111.105p 0.549932mV 925121.251p 0.551813mV 925132.932p 0.5537mV 926026.618p 0.556475mV 926028.765p 0.556475mV 926051.129p 0.558727mV 926075.029p 0.556291mV 926106.136p 0.553674mV 926117.314p 0.554281mV 926125.456p 0.553438mV 926132.196p 0.552473mV 926142.095p 0.550187mV 927001.089p 0.547583mV 927002.986p 0.547583mV 927012.783p 0.548004mV 927019.702p 0.548762mV 927022.102p 0.549153mV 927049.334p 0.555862mV 928030.493p 0.559006mV 928032.209p 0.559006mV 929000.114p 0.548632mV 929050.473p 0.53874mV 930004.89p 0.552014mV 930027.582p 0.54857mV 930058.988p 0.543298mV 930065.803p 0.542977mV 930087.342p 0.543015mV 931009.992p 0.551666mV 931015.295p 0.55122mV 932033.749p 0.557605mV 932048.863p 0.55954mV 932049.229p 0.55954mV 933010.875p 0.549789mV 933021.643p 0.551798mV 933024.472p 0.551798mV 933040.231p 0.558034mV 933040.878p 0.558034mV 934001.13p 0.547446mV 934032.723p 0.549446mV 935010.753p 0.552608mV 935024.694p 0.553139mV 935109.036p 0.564164mV 936001.888p 0.547732mV 936018.062p 0.547842mV 936028.997p 0.548035mV 936050.518p 0.546502mV 936065.331p 0.545137mV 936073.086p 0.54468mV 936086.816p 0.544029mV 936098.879p 0.544194mV 936118.65p 0.543036mV 936131.854p 0.54488mV 936163.347p 0.552514mV 936164.604p 0.552514mV 936174.893p 0.553339mV 936191.178p 0.557169mV 936201.618p 0.558711mV 936241.214p 0.564102mV 936273.955p 0.566432mV 936311.601p 0.5767mV 936319.281p 0.5787mV 936387.796p 0.601578mV 936392.075p 0.603884mV 936417.817p 0.615718mV 936424.82p 0.618mV 936433.387p 0.623646mV 936444.527p 0.629275mV 936451.427p 0.635617mV 936464.218p 0.642673mV 937020.605p 0.547792mV 937023.512p 0.547792mV 938007.52p 0.546596mV 938014.744p 0.546894mV 938023.607p 0.548587mV 938045.564p 0.553385mV 938085.917p 0.555213mV 938171.574p 0.53465mV 939005.365p 0.550133mV 939019.301p 0.550519mV 939025.384p 0.551633mV 939033.766p 0.552737mV 940002.736p 0.550501mV 940004.988p 0.550501mV 940006.06p 0.550574mV 940018.173p 0.549621mV 940029.25p 0.547199mV 940030.392p 0.545437mV 940043.178p 0.543001mV 940044.591p 0.543001mV 941008.496p 0.550591mV 941011.149p 0.551013mV 941014.914p 0.551013mV 941022.687p 0.551488mV 941029.746p 0.552273mV 941040.746p 0.552428mV 941069.484p 0.548283mV 942014.851p 0.547503mV 942019.169p 0.547471mV 942025.954p 0.54631mV 942048.768p 0.539603mV 942053.108p 0.537742mV 944011.062p 0.550629mV 944016.722p 0.551396mV 944044.265p 0.558543mV 945027.455p 0.541354mV 946019.768p 0.551681mV 946033.172p 0.551557mV 946050.635p 0.546266mV 946052.385p 0.546266mV 946062.723p 0.543612mV 946073.807p 0.540946mV 947074.893p 0.547862mV 947150.024p 0.553324mV 948001.977p 0.548331mV 948003.6p 0.548331mV 948040.451p 0.541376mV 948044.582p 0.541376mV 948046.479p 0.54059mV 949041.703p 0.544497mV 949043.842p 0.544497mV 949054.245p 0.544188mV 950005.743p 0.5538mV 950027.548p 0.556238mV 950058.505p 0.561379mV 950077.831p 0.566067mV 951002.79p 0.552115mV 951019.767p 0.551679mV 951029.291p 0.551262mV 951045.606p 0.55261mV 951080.768p 0.559707mV 951113.23p 0.567264mV 952011.533p 0.547827mV 952019.902p 0.547842mV 952020.978p 0.547491mV 952034.293p 0.54569mV 952102.694p 0.543064mV 952113.439p 0.544823mV 952123.27p 0.548028mV 952134.557p 0.550489mV 952139.244p 0.551898mV 952156.38p 0.558974mV 952163.156p 0.560007mV 952183.148p 0.564127mV 952188.979p 0.565519mV 952214.916p 0.577219mV 952222.878p 0.581825mV 952235.421p 0.589296mV 952242.026p 0.59106mV 952268.534p 0.596654mV 952275.413p 0.597679mV 952277.051p 0.597679mV 952277.448p 0.597679mV 952301.739p 0.600134mV 953005.121p 0.551733mV 953007.894p 0.551733mV 953012.101p 0.55129mV 953034.69p 0.553177mV 953062.578p 0.560426mV 954008.681p 0.552769mV 954037.293p 0.552855mV 954037.359p 0.552855mV 954046.797p 0.555554mV 954057.481p 0.557517mV 954091.345p 0.566054mV 954092.534p 0.566054mV 954097.153p 0.566864mV 955001.365p 0.554251mV 955053.97p 0.557646mV 955074.06p 0.561816mV 955079.566p 0.563231mV 956006.533p 0.553386mV 956008.288p 0.553386mV 956043.587p 0.551792mV 956065.095p 0.552936mV 956066.946p 0.552936mV 956105.857p 0.555018mV 956140.347p 0.562853mV 956152.062p 0.5663mV 957037.561p 0.542157mV 957050.07p 0.536907mV 958019.329p 0.548031mV 958026.684p 0.547535mV 958052.676p 0.545389mV 958086.0p 0.537991mV 958091.821p 0.536825mV 959013.39p 0.5508mV 959044.578p 0.54876mV 959047.303p 0.548117mV 959064.662p 0.547648mV 959085.83p 0.54515mV 959096.706p 0.544949mV 959116.565p 0.543062mV 959117.77p 0.543062mV 959146.706p 0.540154mV 960025.364p 0.55265mV 960040.241p 0.55263mV 960040.758p 0.55263mV 960122.842p 0.559046mV 960153.432p 0.553535mV 960158.26p 0.552798mV 960189.299p 0.55309mV 960231.961p 0.55321mV 960235.32p 0.551711mV 960239.667p 0.551711mV 961005.846p 0.552121mV 961059.426p 0.547388mV 962103.22p 0.542519mV 962167.631p 0.562372mV 962169.199p 0.562372mV 962182.907p 0.572254mV 962187.555p 0.575794mV 963030.925p 0.545996mV 963031.983p 0.545996mV 963050.616p 0.548335mV 963061.207p 0.551706mV 963079.06p 0.556596mV 964000.913p 0.550972mV 964038.431p 0.548739mV 964071.835p 0.543856mV 964093.741p 0.544635mV 965000.88p 0.554661mV 965060.231p 0.548681mV 965060.973p 0.548681mV 965071.523p 0.546947mV 965080.351p 0.544473mV 966007.959p 0.550173mV 966076.451p 0.559749mV 966077.266p 0.559749mV 967010.025p 0.55119mV 967047.791p 0.551723mV 967049.148p 0.551723mV 967083.631p 0.553348mV 967092.688p 0.555016mV 967102.495p 0.557418mV 967122.48p 0.561513mV 968019.016p 0.55423mV 968040.828p 0.560014mV 969001.503p 0.547582mV 969006.294p 0.547653mV 969011.132p 0.547358mV 969013.599p 0.547358mV 969016.127p 0.547429mV 969016.34p 0.547429mV 969027.017p 0.546475mV 969037.551p 0.544059mV 969038.791p 0.544059mV 969047.914p 0.541641mV 970000.47p 0.550923mV 970027.95p 0.553375mV 970029.502p 0.553375mV 970040.48p 0.553815mV 970042.216p 0.553815mV 970048.267p 0.554449mV 970060.18p 0.55416mV 970076.479p 0.552046mV 970094.856p 0.548833mV 970108.179p 0.546706mV 970131.071p 0.541404mV 971011.239p 0.547055mV 971011.568p 0.547055mV 971031.943p 0.54542mV 971045.823p 0.544198mV 971065.167p 0.539642mV 972018.422p 0.547634mV 972023.248p 0.548738mV 972027.07p 0.550209mV 972030.159p 0.552046mV 972041.075p 0.556823mV 973017.667p 0.551984mV 973025.927p 0.549315mV 973034.424p 0.54743mV 973057.394p 0.540542mV 974008.584p 0.545896mV 974020.105p 0.548058mV 974020.317p 0.548058mV 974025.401p 0.548778mV 974079.106p 0.555687mV 974084.187p 0.556063mV 974087.122p 0.556809mV 975030.563p 0.556263mV 975031.295p 0.556263mV 975034.951p 0.556263mV 975037.762p 0.556327mV 975069.143p 0.552706mV 975083.625p 0.549252mV 975091.129p 0.546822mV 975109.277p 0.542979mV 976023.643p 0.54714mV 976033.887p 0.545194mV 976047.302p 0.541726mV 976049.6p 0.541726mV 976053.181p 0.539836mV 978016.631p 0.549996mV 978036.869p 0.553589mV 978063.438p 0.561944mV 979012.496p 0.55007mV 979077.357p 0.540652mV 979080.976p 0.539498mV 979097.361p 0.536019mV 979097.714p 0.536019mV 980005.356p 0.553529mV 980031.327p 0.549072mV 980033.682p 0.549072mV 980046.975p 0.544477mV 981047.162p 0.549543mV 981047.66p 0.549543mV 981059.261p 0.552099mV 982023.701p 0.551129mV 982038.545p 0.554353mV 982047.64p 0.556872mV 982051.475p 0.558682mV 982053.005p 0.558682mV 983008.593p 0.554557mV 983023.151p 0.553939mV 983029.518p 0.553974mV 983045.567p 0.55556mV 983055.592p 0.558172mV 983068.044p 0.560782mV 983091.549p 0.573714mV 984007.151p 0.545746mV 984037.713p 0.547711mV 984044.378p 0.548104mV 984073.435p 0.54867mV 984074.289p 0.54867mV 984090.348p 0.548122mV 984091.849p 0.548122mV 984094.552p 0.548122mV 984103.382p 0.549326mV 985003.53p 0.545397mV 985008.802p 0.545454mV 985087.935p 0.533219mV 986008.493p 0.547409mV 986010.051p 0.547037mV 986010.846p 0.547037mV 986038.844p 0.543361mV 986039.265p 0.543361mV 986066.633p 0.537109mV 987015.996p 0.553762mV 987021.74p 0.554052mV 987031.469p 0.553534mV 987093.025p 0.556956mV 987100.851p 0.559349mV 987105.281p 0.56mV 987107.922p 0.56mV 987110.928p 0.561017mV 987136.799p 0.566514mV 988006.337p 0.546453mV 988058.668p 0.556349mV 989016.464p 0.553102mV 989043.627p 0.549396mV 990014.684p 0.548597mV 990029.406p 0.546043mV 990032.477p 0.545679mV 990049.468p 0.543116mV 990079.301p 0.541223mV 990087.986p 0.542273mV 990127.994p 0.545613mV 991006.708p 0.547477mV 991015.102p 0.546504mV 991040.274p 0.539851mV 992006.947p 0.552397mV 992008.788p 0.552397mV 992016.344p 0.551311mV 992032.366p 0.549128mV 992032.866p 0.549128mV 992047.306p 0.545836mV 992074.663p 0.54468mV 993033.688p 0.551521mV 993059.221p 0.554354mV 994007.298p 0.550676mV 994011.15p 0.550981mV 994018.644p 0.551653mV 994037.681p 0.554347mV 994044.492p 0.55539mV 995049.13p 0.559488mV 995063.39p 0.564029mV 996015.289p 0.54807mV 996038.143p 0.547339mV 996084.123p 0.549039mV 996084.241p 0.549039mV 996097.751p 0.545664mV 996100.443p 0.544534mV 996103.935p 0.544534mV 997009.476p 0.548769mV 997009.946p 0.548769mV 997010.736p 0.548377mV 997042.406p 0.548573mV 997086.644p 0.561473mV 998043.791p 0.547818mV 998051.389p 0.544543mV 998073.659p 0.537975mV 999002.328p 0.546362mV 999039.975p 0.546963mV 999064.483p 0.548487mV 999082.918p 0.550489mV)
.ENDS conductors__anyBias-Lk_0_701


.SUBCKT conductors__anyBias-Lk_0_702 bottom out
VrampSppl@0 bottom out pwl(0 0 25.72p 0.563916mV 1001.855p 0.553667mV 1034.061p 0.623876mV 1055.886p 0.641916mV 1057.538p 0.641916mV 2026.505p 0.531548mV 2066.625p 0.566605mV 2122.632p 0.654197mV 3007.185p 0.531811mV 3037.349p 0.496964mV 3049.474p 0.496947mV 3050.894p 0.479355mV 3060.161p 0.444122mV 3072.001p 0.478981mV 4022.201p 0.513182mV 4034.513p 0.513055mV 4035.905p 0.495408mV 4051.896p 0.477482mV 4056.012p 0.459774mV 5042.584p 0.550836mV 5057.084p 0.533435mV 5073.677p 0.480855mV 5088.744p 0.49837mV 5102.911p 0.480591mV 6015.744p 0.570307mV 6016.271p 0.570307mV 6023.999p 0.552737mV 7012.588p 0.518504mV 7023.636p 0.518351mV 7037.055p 0.535581mV 7105.496p 0.533432mV 8010.347p 0.581359mV 8014.016p 0.581359mV 8045.959p 0.5643mV 8079.364p 0.494603mV 8094.871p 0.47719mV 8131.088p 0.441345mV 9039.513p 0.602452mV 9053.145p 0.620286mV 10001.334p 0.54557mV 10003.555p 0.54557mV 10004.789p 0.54557mV 10017.435p 0.493034mV 10042.76p 0.440226mV 11040.322p 0.615797mV 11058.291p 0.633507mV 12012.106p 0.550734mV 12035.263p 0.497767mV 12080.836p 0.548902mV 12092.142p 0.513413mV 13045.803p 0.528801mV 13084.226p 0.545566mV 13101.948p 0.509727mV 14020.248p 0.545618mV 14042.395p 0.510303mV 14058.315p 0.492515mV 14073.732p 0.50968mV 14092.724p 0.543987mV 14097.947p 0.561277mV 15053.084p 0.547718mV 15056.716p 0.530054mV 15063.858p 0.512388mV 15068.717p 0.494717mV 15081.927p 0.476718mV 16003.478p 0.546277mV 16028.766p 0.528983mV 16042.092p 0.476505mV 16056.788p 0.458967mV 16101.273p 0.510211mV 17000.996p 0.548684mV 17001.053p 0.548684mV 17018.193p 0.566412mV 17036.048p 0.566701mV 17036.946p 0.566701mV 17043.945p 0.584354mV 18014.523p 0.514043mV 18021.839p 0.514016mV 18024.116p 0.514016mV 18055.605p 0.56596mV 18088.013p 0.529874mV 19000.708p 0.546879mV 19049.433p 0.494331mV 19076.956p 0.493869mV 19084.825p 0.476194mV 19089.103p 0.45851mV 19091.773p 0.475882mV 20034.417p 0.516214mV 20044.843p 0.516013mV 20059.008p 0.498026mV 21003.46p 0.546885mV 21053.228p 0.582086mV 21068.692p 0.599707mV 21079.404p 0.634974mV 21079.94p 0.634974mV 21080.892p 0.652629mV 22004.729p 0.552726mV 22009.922p 0.535177mV 22010.527p 0.517628mV 22015.692p 0.535194mV 22032.047p 0.51759mV 22089.504p 0.569239mV 22095.764p 0.603946mV 22096.613p 0.603946mV 22110.43p 0.656114mV 22111.787p 0.656114mV 22119.404p 0.638462mV 22120.959p 0.65594mV 22136.846p 0.708558mV 22139.924p 0.708558mV 23053.777p 0.516203mV 23071.079p 0.516141mV 24002.588p 0.547536mV 24009.408p 0.565139mV 24011.078p 0.582743mV 24018.17p 0.600354mV 24022.757p 0.617977mV 24030.299p 0.653269mV 24031.69p 0.653269mV 25013.949p 0.551624mV 25053.03p 0.586951mV 25081.809p 0.552151mV 25091.494p 0.517175mV 25092.102p 0.517175mV 25092.524p 0.517175mV 25092.778p 0.517175mV 25154.966p 0.446666mV 26008.321p 0.564933mV 26010.849p 0.582478mV 26022.684p 0.582479mV 26030.402p 0.54744mV 26033.423p 0.54744mV 26123.972p 0.58421mV 27022.801p 0.583719mV 27034.175p 0.583738mV 28024.551p 0.550897mV 28055.998p 0.638589mV 28077.645p 0.674014mV 28079.498p 0.674014mV 29015.958p 0.568997mV 29035.236p 0.639182mV 29053.438p 0.65694mV 29056.505p 0.674607mV 30020.296p 0.586546mV 30032.193p 0.586529mV 30070.331p 0.586993mV 30072.591p 0.586993mV 30080.476p 0.552142mV 30088.4p 0.53474mV 30125.906p 0.465267mV 30130.272p 0.482804mV 30138.477p 0.465195mV 30152.183p 0.44736mV 31042.162p 0.553777mV 31044.957p 0.553777mV 31056.393p 0.571305mV 31072.539p 0.623957mV 31118.294p 0.607241mV 32004.293p 0.545789mV 32036.269p 0.528585mV 32040.048p 0.546181mV 32076.305p 0.49355mV 32087.593p 0.493374mV 33033.707p 0.546488mV 33037.616p 0.56407mV 33109.521p 0.458782mV 33110.208p 0.4411mV 33111.174p 0.4411mV 33116.738p 0.423414mV 34023.371p 0.55029mV 34034.611p 0.515306mV 34041.457p 0.550532mV 34101.445p 0.586228mV 34134.895p 0.552175mV 34144.526p 0.517583mV 34188.892p 0.431753mV 34204.941p 0.449601mV 34206.608p 0.432105mV 34228.866p 0.432162mV 35010.318p 0.584942mV 35027.133p 0.567416mV 35068.016p 0.56826mV 35083.132p 0.551379mV 36012.443p 0.518433mV 36028.421p 0.500934mV 36034.351p 0.483363mV 36040.845p 0.518397mV 36044.604p 0.518397mV 36045.654p 0.535875mV 36047.357p 0.535875mV 36101.901p 0.551651mV 37034.503p 0.519044mV 37064.518p 0.483726mV 37064.967p 0.483726mV 37069.758p 0.501172mV 38018.047p 0.501559mV 38024.148p 0.519153mV 38062.01p 0.518894mV 38090.622p 0.483079mV 39001.841p 0.551474mV 39012.658p 0.551421mV 39062.742p 0.586127mV 39076.946p 0.603677mV 40016.2p 0.563122mV 40024.749p 0.580635mV 40033.195p 0.580574mV 40064.08p 0.545434mV 40086.767p 0.598075mV 40135.86p 0.528624mV 40192.8p 0.511824mV 40199.67p 0.52937mV 40223.348p 0.511651mV 40227.777p 0.529147mV 41013.633p 0.518621mV 41031.308p 0.588676mV 41044.881p 0.58859mV 41064.623p 0.553379mV 42012.041p 0.515678mV 42015.364p 0.49805mV 42025.474p 0.497859mV 42032.611p 0.515283mV 42051.119p 0.51456mV 43015.387p 0.568541mV 43026.046p 0.533532mV 43036.974p 0.568761mV 43050.841p 0.586514mV 43058.013p 0.569047mV 43070.057p 0.551846mV 43093.536p 0.552459mV 43094.774p 0.552459mV 43099.332p 0.53512mV 43116.991p 0.500872mV 43124.077p 0.483538mV 43126.26p 0.501259mV 43143.183p 0.484242mV 43184.899p 0.415001mV 43185.127p 0.397465mV 43191.275p 0.415023mV 44001.572p 0.552018mV 44022.652p 0.481749mV 44028.25p 0.499268mV 44039.859p 0.499105mV 45060.654p 0.620411mV 46018.625p 0.532493mV 46021.475p 0.514938mV 46043.934p 0.514874mV 46050.657p 0.514799mV 46068.025p 0.497003mV 46069.819p 0.497003mV 47028.716p 0.566511mV 47037.288p 0.566577mV 47059.702p 0.531704mV 47079.489p 0.531904mV 47116.969p 0.531603mV 49009.211p 0.531673mV 49045.618p 0.56735mV 49078.985p 0.568117mV 50017.494p 0.534662mV 50026.67p 0.569804mV 50043.275p 0.587405mV 50056.082p 0.569959mV 50067.009p 0.534985mV 50123.799p 0.447874mV 50127.21p 0.465406mV 50177.958p 0.568867mV 50180.33p 0.58612mV 51007.469p 0.571068mV 51008.774p 0.571068mV 51054.096p 0.519mV 51062.386p 0.519095mV 51082.781p 0.519174mV 51095.646p 0.501519mV 51098.141p 0.501519mV 51100.173p 0.519035mV 51135.134p 0.535967mV 51140.661p 0.553384mV 51144.257p 0.553384mV 51151.516p 0.55311mV 51153.113p 0.55311mV 51153.908p 0.55311mV 51158.664p 0.535432mV 54018.465p 0.532485mV 54066.007p 0.461766mV 55008.393p 0.570595mV 55028.838p 0.605881mV 55030.66p 0.588426mV 55042.162p 0.588691mV 55044.217p 0.588691mV 55044.573p 0.588691mV 55058.227p 0.606765mV 56025.342p 0.564939mV 56049.085p 0.565031mV 56067.199p 0.565295mV 56073.911p 0.547839mV 56083.391p 0.548053mV 56091.45p 0.548263mV 56118.059p 0.566505mV 56126.596p 0.601927mV 56127.243p 0.601927mV 57015.75p 0.493147mV 57059.358p 0.527344mV 58001.922p 0.547253mV 58032.958p 0.582276mV 58073.632p 0.54746mV 58087.178p 0.565189mV 58149.34p 0.56701mV 59004.664p 0.553746mV 59026.732p 0.57136mV 59075.93p 0.607324mV 59076.075p 0.607324mV 60049.539p 0.563202mV 60068.255p 0.528226mV 60068.712p 0.528226mV 60072.656p 0.545816mV 60107.499p 0.45792mV 60111.252p 0.440267mV 61027.455p 0.535538mV 61032.435p 0.553038mV 61037.351p 0.535413mV 61042.273p 0.517787mV 61062.414p 0.587612mV 61080.252p 0.587229mV 61087.948p 0.604714mV 61090.359p 0.622209mV 61108.138p 0.604561mV 61136.17p 0.604715mV 61150.751p 0.587346mV 61161.837p 0.552389mV 61165.235p 0.570027mV 61179.945p 0.570184mV 61195.143p 0.570476mV 61206.291p 0.570601mV 61213.497p 0.588222mV 61213.928p 0.588222mV 61219.863p 0.605848mV 61230.463p 0.623698mV 61232.883p 0.623698mV 61237.827p 0.606297mV 62003.562p 0.549906mV 62011.93p 0.514841mV 62037.787p 0.5324mV 62045.233p 0.532359mV 62087.319p 0.531646mV 62126.501p 0.565375mV 63012.319p 0.548911mV 63013.531p 0.548911mV 63020.906p 0.584044mV 63028.41p 0.566497mV 63059.177p 0.531568mV 63062.592p 0.549155mV 63063.147p 0.549155mV 63099.378p 0.531763mV 63115.196p 0.602123mV 63132.153p 0.584794mV 63136.414p 0.602465mV 64006.58p 0.563619mV 64057.102p 0.634349mV 65015.784p 0.566034mV 65028.269p 0.601221mV 65052.928p 0.689415mV 66023.591p 0.622594mV 66023.997p 0.622594mV 66033.397p 0.587525mV 66039.661p 0.605145mV 66102.701p 0.589481mV 67013.246p 0.584321mV 67017.825p 0.601933mV 67032.168p 0.584634mV 67046.416p 0.637648mV 67051.152p 0.655335mV 68028.29p 0.600487mV 68050.301p 0.583512mV 68058.13p 0.601225mV 69003.892p 0.550741mV 69015.323p 0.568098mV 69015.928p 0.568098mV 69033.712p 0.550329mV 69038.269p 0.56782mV 69039.736p 0.56782mV 69069.756p 0.60252mV 69077.268p 0.637535mV 69088.667p 0.637525mV 69119.377p 0.603037mV 69127.166p 0.603404mV 70016.651p 0.532315mV 70051.576p 0.514203mV 70057.474p 0.496522mV 70062.069p 0.478834mV 71021.11p 0.583545mV 71045.94p 0.636345mV 71046.486p 0.636345mV 71053.554p 0.653978mV 71064.75p 0.654216mV 72032.788p 0.519323mV 72040.341p 0.55448mV 72059.701p 0.53694mV 72087.006p 0.466541mV 72108.235p 0.465971mV 73008.653p 0.569776mV 73019.628p 0.534727mV 73034.642p 0.552386mV 73044.473p 0.587581mV 73059.929p 0.570213mV 73081.588p 0.553236mV 73104.804p 0.518664mV 73171.191p 0.519399mV 73184.735p 0.519353mV 73188.879p 0.50176mV 73197.064p 0.501683mV 73198.898p 0.501683mV 74010.65p 0.549976mV 74046.097p 0.637981mV 74065.744p 0.638467mV 75005.045p 0.569556mV 75012.536p 0.55202mV 75015.257p 0.569612mV 75039.104p 0.569774mV 75041.091p 0.552265mV 75047.93p 0.534766mV 75052.595p 0.552384mV 75058.254p 0.534881mV 75059.427p 0.534881mV 75063.036p 0.517381mV 75067.605p 0.534992mV 75082.475p 0.587791mV 75102.239p 0.552968mV 75107.835p 0.535517mV 75111.727p 0.518073mV 75119.734p 0.535732mV 75128.107p 0.535933mV 75147.485p 0.501235mV 75211.223p 0.448064mV 76003.46p 0.550574mV 76014.423p 0.51535mV 76014.443p 0.51535mV 76018.068p 0.53285mV 76055.663p 0.602675mV 76084.306p 0.55038mV 76085.355p 0.532921mV 76086.878p 0.532921mV 76103.342p 0.51562mV 76111.755p 0.550832mV 76140.177p 0.515839mV 76145.269p 0.533373mV 76149.221p 0.533373mV 76164.267p 0.550814mV 76164.544p 0.550814mV 76179.898p 0.568306mV 76187.221p 0.533168mV 76199.732p 0.568282mV 76202.042p 0.550717mV 76247.007p 0.462634mV 77000.528p 0.546862mV 77069.526p 0.599443mV 77092.787p 0.582662mV 78022.715p 0.553425mV 78046.418p 0.500228mV 79000.5p 0.554429mV 79011.95p 0.554305mV 79031.15p 0.554033mV 79031.835p 0.554033mV 79069.581p 0.535917mV 80012.981p 0.513381mV 80013.538p 0.513381mV 80064.133p 0.443099mV 81005.589p 0.534062mV 81060.326p 0.517059mV 81077.823p 0.534769mV 81111.558p 0.55262mV 81158.182p 0.535449mV 81168.376p 0.535538mV 81171.442p 0.518017mV 81181.389p 0.482972mV 81202.113p 0.482968mV 81235.019p 0.535044mV 81245.394p 0.534793mV 81278.492p 0.533814mV 82077.368p 0.53363mV 82091.648p 0.550905mV 82107.767p 0.568074mV 82116.145p 0.602863mV 82122.216p 0.585175mV 82131.769p 0.620002mV 82138.117p 0.637429mV 82141.907p 0.654878mV 82141.945p 0.654878mV 82207.784p 0.672488mV 82207.927p 0.672488mV 82229.14p 0.60287mV 83017.574p 0.600741mV 83059.922p 0.601343mV 83061.966p 0.583957mV 84015.001p 0.563842mV 84044.429p 0.616619mV 84070.149p 0.547445mV 84079.704p 0.565202mV 85003.324p 0.553135mV 85018.368p 0.535578mV 85068.0p 0.605915mV 85082.6p 0.553469mV 85090.57p 0.588785mV 85128.095p 0.572436mV 86020.292p 0.514762mV 86021.514p 0.514762mV 87049.365p 0.496443mV 87067.516p 0.460841mV 88009.228p 0.563302mV 88044.25p 0.511229mV 88113.05p 0.547225mV 88115.659p 0.529764mV 88115.723p 0.529764mV 88151.696p 0.407444mV 90002.235p 0.551285mV 90036.927p 0.56851mV 90049.821p 0.533299mV 90099.843p 0.602979mV 90100.834p 0.58545mV 90101.026p 0.58545mV 90106.666p 0.603058mV 90109.809p 0.603058mV 90113.985p 0.585557mV 91014.057p 0.587406mV 91031.931p 0.587469mV 91048.596p 0.570092mV 91086.103p 0.46541mV 91108.847p 0.465206mV 91117.218p 0.464942mV 92026.784p 0.603576mV 92031.955p 0.621159mV 92045.834p 0.638922mV 92050.158p 0.656588mV 93001.243p 0.549144mV 93065.019p 0.567688mV 93088.461p 0.568393mV 93089.304p 0.568393mV 93095.601p 0.568792mV 94020.845p 0.582108mV 94048.223p 0.600066mV 94080.801p 0.548676mV 94081.689p 0.548676mV 94173.866p 0.517568mV 94177.3p 0.535291mV 94184.447p 0.553016mV 95024.149p 0.513872mV 95044.605p 0.478578mV 96003.3p 0.553021mV 96014.274p 0.517793mV 96034.514p 0.517424mV 96035.949p 0.534813mV 97050.87p 0.587243mV 97050.942p 0.587243mV 97054.944p 0.587243mV 97100.899p 0.552915mV 97106.483p 0.535436mV 97123.924p 0.553225mV 97158.028p 0.606516mV 97162.639p 0.624199mV 98031.581p 0.483188mV 99007.224p 0.530357mV 99052.423p 0.442269mV 100006.277p 0.530925mV 100017.402p 0.495852mV 100020.116p 0.478296mV 100034.969p 0.513354mV 100059.74p 0.495323mV 101022.207p 0.550976mV 101024.436p 0.550976mV 101043.774p 0.586153mV 101047.288p 0.603751mV 101047.662p 0.603751mV 101067.894p 0.604076mV 101084.801p 0.551968mV 101097.47p 0.535077mV 101112.527p 0.518233mV 101120.804p 0.518667mV 101131.635p 0.55416mV 102002.314p 0.546731mV 102027.307p 0.564104mV 102039.251p 0.56406mV 102065.533p 0.634432mV 102080.867p 0.582132mV 103008.859p 0.53035mV 103018.491p 0.49521mV 103021.571p 0.477624mV 103023.332p 0.477624mV 104014.603p 0.545633mV 104016.213p 0.528134mV 104031.985p 0.510718mV 104059.665p 0.563396mV 104072.527p 0.545797mV 104131.922p 0.545968mV 104153.832p 0.510946mV 104153.843p 0.510946mV 104214.055p 0.545581mV 104232.879p 0.545279mV 104279.113p 0.526589mV 104290.695p 0.578419mV 104307.336p 0.595158mV 104353.244p 0.645555mV 104355.319p 0.627801mV 104359.461p 0.627801mV 105006.172p 0.56429mV 105033.043p 0.546846mV 105036.056p 0.529316mV 105066.362p 0.529315mV 105069.468p 0.529315mV 105071.185p 0.54683mV 105100.464p 0.581712mV 105120.373p 0.652009mV 105139.84p 0.704924mV 107008.504p 0.570684mV 107037.971p 0.570658mV 107038.576p 0.570658mV 107055.907p 0.570958mV 107080.663p 0.553876mV 107086.704p 0.571538mV 107098.848p 0.536683mV 107145.099p 0.502861mV 107205.596p 0.502594mV 108004.742p 0.552988mV 108015.985p 0.535331mV 110027.153p 0.599213mV 110030.986p 0.58169mV 110065.503p 0.564727mV 110082.137p 0.547493mV 111012.171p 0.581421mV 111021.434p 0.581421mV 111040.913p 0.546418mV 111062.796p 0.546598mV 111064.856p 0.546598mV 111064.993p 0.546598mV 111075.377p 0.599355mV 112033.015p 0.58792mV 112040.344p 0.623125mV 112050.08p 0.62329mV 112065.671p 0.57112mV 113011.879p 0.546901mV 113019.12p 0.529317mV 113075.791p 0.634412mV 113080.461p 0.652035mV 113085.233p 0.669676mV 113088.183p 0.669676mV 113091.056p 0.68733mV 113097.002p 0.669928mV 114021.373p 0.5523mV 114037.777p 0.570003mV 114049.2p 0.570153mV 114054.199p 0.552697mV 114062.827p 0.517817mV 114066.421p 0.500374mV 114091.598p 0.518293mV 114097.721p 0.535904mV 114115.499p 0.465824mV 114159.532p 0.43016mV 115016.919p 0.528275mV 115027.964p 0.528129mV 115028.814p 0.528129mV 115036.481p 0.563071mV 115044.328p 0.580534mV 115048.493p 0.562892mV 115052.151p 0.545259mV 115085.989p 0.491784mV 115089.317p 0.491784mV 116014.759p 0.554097mV 116042.188p 0.519008mV 116114.439p 0.587308mV 116118.883p 0.569581mV 116121.625p 0.551857mV 116129.969p 0.569191mV 116130.13p 0.586504mV 117000.759p 0.55339mV 118003.334p 0.548216mV 118058.711p 0.4602mV 119082.697p 0.589041mV 119082.925p 0.589041mV 119090.504p 0.58938mV 120034.783p 0.514918mV 120043.228p 0.479637mV 120044.583p 0.479637mV 121000.335p 0.547097mV 121001.428p 0.547097mV 121014.222p 0.582236mV 121015.926p 0.599813mV 121024.435p 0.582282mV 121033.39p 0.617515mV 121034.281p 0.617515mV 121038.527p 0.600044mV 121042.732p 0.582609mV 121055.717p 0.600611mV 121055.901p 0.600611mV 122037.675p 0.6069mV 123011.204p 0.551352mV 123030.731p 0.586624mV 123034.119p 0.586624mV 123054.462p 0.657183mV 124014.425p 0.511793mV 124041.141p 0.51152mV 124067.661p 0.493168mV 125024.224p 0.6198mV 125066.288p 0.567944mV 125081.682p 0.62099mV 126005.892p 0.564607mV 126043.885p 0.547039mV 126066.462p 0.599791mV 126075.304p 0.599904mV 126104.464p 0.583089mV 127008.915p 0.528006mV 127010.063p 0.51043mV 127026.938p 0.492759mV 127046.949p 0.492314mV 127052.617p 0.509682mV 128005.293p 0.53307mV 128025.119p 0.497901mV 128030.473p 0.48029mV 128030.94p 0.48029mV 128037.969p 0.462664mV 129004.638p 0.553206mV 129031.481p 0.588566mV 129037.411p 0.606169mV 129048.428p 0.641415mV 129056.957p 0.606554mV 129059.314p 0.606554mV 130002.329p 0.546257mV 130003.542p 0.546257mV 130052.521p 0.545678mV 130054.629p 0.545678mV 130056.96p 0.563186mV 130063.131p 0.58069mV 130069.501p 0.5982mV 130070.947p 0.580603mV 130074.8p 0.580603mV 130113.856p 0.545688mV 130131.661p 0.510846mV 130146.807p 0.493406mV 130151.24p 0.475835mV 130158.997p 0.458245mV 130165.645p 0.458106mV 131004.275p 0.546413mV 131005.085p 0.563966mV 131029.625p 0.528825mV 131058.595p 0.598792mV 131087.835p 0.528631mV 131091.941p 0.546236mV 131130.725p 0.581933mV 131133.957p 0.581933mV 132013.836p 0.553054mV 132058.222p 0.571108mV 132072.893p 0.55389mV 132083.855p 0.554151mV 132095.079p 0.501971mV 132115.148p 0.502485mV 132117.348p 0.502485mV 132151.21p 0.48556mV 132171.527p 0.48578mV 132208.058p 0.50333mV 132250.612p 0.414975mV 133002.2p 0.554321mV 133009.079p 0.536773mV 133012.235p 0.519226mV 133023.823p 0.484102mV 133028.954p 0.466514mV 133041.531p 0.448715mV 133042.919p 0.448715mV 134042.404p 0.616655mV 134056.607p 0.564313mV 134060.96p 0.582003mV 134082.286p 0.547623mV 135005.476p 0.563302mV 135046.958p 0.598109mV 135053.743p 0.615675mV 135066.058p 0.633382mV 135066.471p 0.633382mV 136099.244p 0.464194mV 136114.283p 0.446312mV 136116.85p 0.463699mV 136123.98p 0.445984mV 137046.888p 0.533098mV 137047.287p 0.533098mV 137077.421p 0.532903mV 137098.637p 0.497462mV 137118.723p 0.496915mV 138034.696p 0.58302mV 138061.369p 0.548087mV 138063.801p 0.548087mV 138076.44p 0.565896mV 138090.331p 0.513597mV 138107.021p 0.496368mV 138131.794p 0.514169mV 138137.146p 0.531761mV 138141.525p 0.549347mV 138163.687p 0.549543mV 138171.329p 0.549743mV 138193.827p 0.585356mV 138202.767p 0.585751mV 139000.184p 0.551674mV 139052.382p 0.552262mV 139067.604p 0.534785mV 139076.465p 0.569963mV 139086.389p 0.605154mV 139100.812p 0.587844mV 139100.963p 0.587844mV 140018.016p 0.528314mV 140032.152p 0.58093mV 140037.726p 0.598473mV 140059.892p 0.633685mV 140067.757p 0.668956mV 141020.724p 0.515455mV 141046.101p 0.567749mV 141069.515p 0.567372mV 141096.61p 0.60203mV 141097.245p 0.60203mV 141122.162p 0.584438mV 141126.18p 0.566866mV 141128.231p 0.566866mV 141155.813p 0.56674mV 141204.98p 0.618855mV 141226.03p 0.671447mV 142004.13p 0.549672mV 142041.567p 0.514215mV 142058.877p 0.496327mV 143028.423p 0.497756mV 144050.579p 0.554153mV 144094.019p 0.553565mV 144126.177p 0.535121mV 145003.451p 0.551941mV 145005.313p 0.569524mV 145038.813p 0.640072mV 145056.267p 0.605646mV 146013.876p 0.553133mV 146034.465p 0.553369mV 146035.379p 0.535848mV 146036.505p 0.535848mV 146061.194p 0.553527mV 146064.195p 0.553527mV 146101.794p 0.588892mV 146121.75p 0.589447mV 147018.091p 0.569202mV 147018.277p 0.569202mV 147031.942p 0.516703mV 147037.339p 0.534315mV 147039.009p 0.534315mV 147057.713p 0.53441mV 148009.069p 0.529697mV 148030.958p 0.511896mV 149016.102p 0.566148mV 149019.626p 0.566148mV 149024.873p 0.58365mV 149027.874p 0.566043mV 149034.0p 0.583569mV 149047.571p 0.6011mV 149058.522p 0.601193mV 149073.781p 0.583955mV 149074.213p 0.583955mV 149104.622p 0.54999mV 150021.94p 0.554418mV 150050.797p 0.589713mV 150080.114p 0.590335mV 151007.13p 0.564926mV 151048.242p 0.600766mV 151058.834p 0.636135mV 152008.192p 0.536186mV 152008.981p 0.536186mV 152012.124p 0.553686mV 152043.865p 0.658773mV 152044.905p 0.658773mV 152045.841p 0.676361mV 152059.499p 0.711605mV 152060.646p 0.69417mV 153001.316p 0.552636mV 153008.555p 0.570228mV 153010.799p 0.587819mV 153013.512p 0.587819mV 153052.04p 0.588754mV 154050.299p 0.549681mV 154098.208p 0.531417mV 154127.32p 0.49544mV 155003.167p 0.552634mV 155005.652p 0.535034mV 155026.262p 0.534853mV 155031.703p 0.55236mV 155037.163p 0.534742mV 155063.179p 0.516776mV 155074.221p 0.481434mV 155083.082p 0.446061mV 156006.405p 0.531729mV 156007.571p 0.531729mV 156028.49p 0.566683mV 156034.384p 0.584188mV 156035.101p 0.601699mV 156036.091p 0.601699mV 156044.839p 0.619225mV 156079.735p 0.602027mV 156086.222p 0.602332mV 156094.963p 0.584974mV 156098.061p 0.602702mV 157007.514p 0.533559mV 157022.668p 0.515888mV 158000.348p 0.548822mV 158017.646p 0.495956mV 159017.883p 0.602953mV 159029.115p 0.567999mV 159048.905p 0.638679mV 160043.143p 0.514446mV 160071.139p 0.548984mV 160097.597p 0.495623mV 160108.172p 0.495253mV 161003.009p 0.546348mV 161009.122p 0.563872mV 161020.181p 0.54624mV 161029.242p 0.528677mV 161063.288p 0.546183mV 161145.772p 0.598594mV 161159.152p 0.56372mV 162011.805p 0.554334mV 162023.649p 0.554295mV 162042.885p 0.554279mV 162056.266p 0.571903mV 163019.815p 0.528994mV 163023.445p 0.546526mV 163032.641p 0.546455mV 163056.444p 0.563931mV 163063.909p 0.58149mV 163102.473p 0.652183mV 164009.625p 0.569233mV 164056.807p 0.605473mV 164061.578p 0.588147mV 165008.409p 0.56949mV 165015.548p 0.569506mV 165036.916p 0.604813mV 165046.32p 0.605013mV 165059.639p 0.640368mV 166017.263p 0.49863mV 166018.195p 0.49863mV 166041.715p 0.480477mV 167017.084p 0.498293mV 167020.507p 0.480701mV 168016.912p 0.603486mV 168020.94p 0.585959mV 168049.479p 0.568862mV 168062.044p 0.586852mV 168069.295p 0.60456mV 168073.944p 0.622272mV 168074.594p 0.622272mV 169003.612p 0.54887mV 169030.529p 0.583857mV 169054.477p 0.584053mV 169081.195p 0.584535mV 169105.768p 0.567652mV 169105.989p 0.567652mV 169107.356p 0.567652mV 169107.82p 0.567652mV 169123.53p 0.550684mV 169126.608p 0.533358mV 169129.541p 0.533358mV 169134.416p 0.551098mV 170034.506p 0.580389mV 170044.807p 0.61546mV 170067.545p 0.633265mV 171000.861p 0.545874mV 171011.225p 0.581059mV 171024.716p 0.616271mV 171030.998p 0.616441mV 172014.259p 0.54614mV 172019.881p 0.563725mV 172028.085p 0.563784mV 172044.392p 0.581468mV 172059.687p 0.529008mV 172074.627p 0.58193mV 172075.767p 0.599579mV 173023.125p 0.516387mV 173063.693p 0.621953mV 174026.348p 0.537093mV 174048.624p 0.537231mV 174067.444p 0.572485mV 174073.465p 0.590103mV 174088.043p 0.572806mV 174089.314p 0.572806mV 174090.838p 0.555378mV 174126.389p 0.504013mV 174130.399p 0.521746mV 174141.216p 0.48709mV 174153.367p 0.487466mV 174186.754p 0.541344mV 174208.838p 0.472197mV 175031.318p 0.589286mV 175035.635p 0.571838mV 175036.688p 0.571838mV 175049.915p 0.607184mV 176025.587p 0.499745mV 176029.013p 0.499745mV 176052.298p 0.516864mV 176066.844p 0.498861mV 177056.699p 0.636808mV 177059.016p 0.636808mV 178009.82p 0.535766mV 178046.641p 0.64159mV 179029.495p 0.49439mV 179043.27p 0.441455mV 179044.949p 0.441455mV 180006.238p 0.571733mV 180008.594p 0.571733mV 180036.525p 0.536385mV 180043.831p 0.553904mV 180066.983p 0.536002mV 180098.843p 0.535224mV 181001.239p 0.550756mV 181004.96p 0.550756mV 181015.785p 0.568234mV 181030.881p 0.585746mV 181086.106p 0.498697mV 181116.361p 0.499012mV 181129.065p 0.463897mV 181140.874p 0.446188mV 182004.632p 0.553885mV 182027.558p 0.501039mV 183040.85p 0.549748mV 183051.645p 0.549728mV 183077.864p 0.496898mV 183079.024p 0.496898mV 183113.808p 0.583905mV 183118.309p 0.601314mV 183129.37p 0.636171mV 183134.489p 0.618527mV 183140.14p 0.653529mV 183163.915p 0.618478mV 183189.124p 0.671694mV 184009.203p 0.56658mV 184015.701p 0.531573mV 184030.773p 0.549292mV 184076.362p 0.531846mV 184077.354p 0.531846mV 184083.523p 0.549377mV 184113.729p 0.549184mV 184152.444p 0.619363mV 184171.994p 0.689963mV 185000.97p 0.545852mV 185009.01p 0.563412mV 185017.809p 0.563419mV 185021.511p 0.545883mV 185039.269p 0.56354mV 185063.356p 0.581401mV 185075.383p 0.599312mV 186028.332p 0.570982mV 186036.027p 0.606025mV 186040.934p 0.623565mV 186070.599p 0.659096mV 186075.755p 0.641728mV 186076.243p 0.641728mV 187009.29p 0.536384mV 187020.207p 0.518913mV 187037.366p 0.501341mV 187064.839p 0.448307mV 188001.609p 0.55074mV 188040.497p 0.621614mV 189060.202p 0.657979mV 189062.209p 0.657979mV 190005.682p 0.569848mV 190044.406p 0.587064mV 190066.039p 0.569348mV 190073.008p 0.551767mV 190136.443p 0.498495mV 190148.092p 0.498165mV 190153.415p 0.515491mV 191013.555p 0.582626mV 192006.32p 0.568884mV 192010.582p 0.551384mV 192026.589p 0.534039mV 192034.259p 0.551674mV 192064.473p 0.552263mV 192117.43p 0.571479mV 193054.729p 0.620994mV 194000.073p 0.552944mV 194043.853p 0.517243mV 194048.718p 0.499538mV 195010.597p 0.513487mV 195046.013p 0.495876mV 196067.053p 0.573151mV 196070.818p 0.555849mV 196078.396p 0.573601mV 197000.188p 0.551497mV 197020.159p 0.551677mV 197039.093p 0.56944mV 197085.802p 0.535626mV 197090.082p 0.553319mV 197102.311p 0.553629mV 198009.032p 0.529206mV 198025.988p 0.494201mV 198033.39p 0.511736mV 198046.973p 0.564224mV 198099.18p 0.528282mV 199038.186p 0.532291mV 199050.304p 0.550007mV 199054.939p 0.550007mV 199088.091p 0.568101mV 199098.669p 0.603436mV 200033.334p 0.585539mV 200044.318p 0.585613mV 200097.438p 0.56969mV 201052.986p 0.51155mV 201055.613p 0.493834mV 202004.684p 0.549655mV 202010.015p 0.549695mV 202011.78p 0.549695mV 202023.229p 0.54972mV 202024.521p 0.54972mV 202041.484p 0.620015mV 202042.814p 0.620015mV 202057.806p 0.567579mV 203025.354p 0.530044mV 203062.359p 0.476687mV 204003.607p 0.550761mV 204003.917p 0.550761mV 205030.381p 0.511242mV 205054.484p 0.476143mV 206003.286p 0.54587mV 206056.292p 0.598509mV 206072.86p 0.581117mV 206092.849p 0.581521mV 206110.137p 0.582189mV 206112.595p 0.582189mV 206119.619p 0.564885mV 207020.452p 0.552825mV 207028.346p 0.53521mV 207040.629p 0.552554mV 207041.961p 0.552554mV 207064.452p 0.517026mV 207081.562p 0.516422mV 208012.325p 0.553481mV 208030.433p 0.553747mV 208046.307p 0.536374mV 208056.643p 0.501382mV 208129.619p 0.535391mV 208134.397p 0.517661mV 208138.864p 0.53498mV 209022.067p 0.552413mV 209031.986p 0.552324mV 209032.53p 0.552324mV 209033.029p 0.552324mV 209037.342p 0.56983mV 209050.081p 0.587246mV 209066.028p 0.569598mV 209093.802p 0.622288mV 209112.805p 0.622736mV 210005.429p 0.566503mV 210069.371p 0.566126mV 210093.155p 0.548727mV 210131.421p 0.584042mV 210132.476p 0.584042mV 210142.53p 0.549073mV 210143.667p 0.549073mV 210147.598p 0.566714mV 210154.111p 0.584354mV 210154.174p 0.584354mV 210188.649p 0.532576mV 210192.46p 0.550266mV 210194.386p 0.550266mV 210200.033p 0.55056mV 210210.778p 0.58595mV 210223.766p 0.586299mV 211055.839p 0.56492mV 211082.048p 0.547727mV 211097.162p 0.530409mV 211113.513p 0.548175mV 211142.35p 0.618934mV 211147.755p 0.601539mV 213023.015p 0.583955mV 213032.877p 0.584112mV 213054.095p 0.549476mV 213065.376p 0.602563mV 214032.931p 0.654549mV 214033.17p 0.654549mV 215002.955p 0.549716mV 215049.704p 0.567443mV 215113.186p 0.51652mV 215124.527p 0.516883mV 216007.708p 0.528895mV 216028.038p 0.529073mV 216028.101p 0.529073mV 216037.193p 0.52912mV 216054.693p 0.546683mV 216060.973p 0.511535mV 216084.349p 0.511364mV 216101.714p 0.510884mV 217056.046p 0.571454mV 217083.794p 0.589454mV 218058.709p 0.461539mV 218076.946p 0.460937mV 218077.464p 0.460937mV 219063.43p 0.589697mV 219078.682p 0.607756mV 219082.237p 0.625483mV 220003.46p 0.552813mV 220026.39p 0.570585mV 220038.344p 0.570706mV 220044.721p 0.553216mV 220064.967p 0.553568mV 220069.036p 0.536127mV 220078.538p 0.536359mV 220079.048p 0.536359mV 220137.554p 0.431149mV 220141.447p 0.413473mV 221048.993p 0.605496mV 221060.443p 0.552903mV 221086.731p 0.535556mV 221106.043p 0.570718mV 221126.046p 0.535739mV 221132.174p 0.518235mV 221133.561p 0.518235mV 221141.602p 0.518321mV 221155.275p 0.535952mV 221187.781p 0.535995mV 221210.424p 0.623942mV 221221.709p 0.624115mV 221228.054p 0.606694mV 221237.613p 0.642095mV 222002.324p 0.545536mV 222009.792p 0.563055mV 222020.306p 0.545381mV 222037.982p 0.527674mV 222076.893p 0.527027mV 223001.016p 0.547891mV 223002.388p 0.547891mV 223011.862p 0.5129mV 223029.266p 0.495459mV 223045.705p 0.530451mV 223052.447p 0.547936mV 223053.899p 0.547936mV 223076.931p 0.63542mV 223100.667p 0.723438mV 224013.676p 0.551082mV 224039.16p 0.568986mV 224068.954p 0.640038mV 225022.958p 0.547292mV 225025.031p 0.564908mV 225063.82p 0.618246mV 225065.161p 0.600887mV 226028.327p 0.532931mV 226069.514p 0.461848mV 227036.448p 0.563005mV 227069.697p 0.527964mV 227069.752p 0.527964mV 227069.785p 0.527964mV 227092.124p 0.580767mV 227106.572p 0.633648mV 228005.539p 0.529199mV 228013.571p 0.546807mV 228037.659p 0.599719mV 228039.241p 0.599719mV 228067.259p 0.600424mV 228071.204p 0.583078mV 228077.688p 0.565773mV 229008.547p 0.569666mV 229009.025p 0.569666mV 229071.388p 0.517607mV 229108.134p 0.500219mV 229152.54p 0.446761mV 229158.856p 0.429076mV 230019.785p 0.564092mV 230027.184p 0.599159mV 230037.357p 0.56404mV 230041.473p 0.546505mV 230052.207p 0.54657mV 230067.687p 0.529117mV 230072.645p 0.546708mV 230085.757p 0.49409mV 230087.367p 0.49409mV 230101.393p 0.511603mV 230121.684p 0.581555mV 230146.493p 0.598973mV 230152.112p 0.616585mV 230152.989p 0.616585mV 230159.549p 0.599099mV 230182.876p 0.582194mV 230183.462p 0.582194mV 230197.789p 0.530091mV 230211.628p 0.548197mV 231007.072p 0.568191mV 231007.555p 0.568191mV 231015.427p 0.532985mV 231032.096p 0.515276mV 231041.766p 0.515091mV 232008.378p 0.565675mV 232014.168p 0.583262mV 232018.62p 0.600856mV 232028.431p 0.600969mV 233018.508p 0.570958mV 233036.481p 0.571048mV 234037.001p 0.57001mV 234045.007p 0.569957mV 234093.843p 0.587418mV 234110.64p 0.587484mV 234114.612p 0.587484mV 234120.229p 0.622702mV 234142.551p 0.623159mV 234143.297p 0.623159mV 235000.622p 0.551048mV 235016.957p 0.568618mV 235028.786p 0.568677mV 235034.765p 0.551168mV 236078.124p 0.564358mV 236091.601p 0.546647mV 236120.365p 0.511167mV 236132.905p 0.475858mV 236137.422p 0.493273mV 236148.76p 0.457867mV 237027.808p 0.532338mV 237043.959p 0.514522mV 237091.141p 0.583332mV 237095.783p 0.600782mV 237126.275p 0.565081mV 237137.359p 0.564821mV 238010.988p 0.551369mV 238017.421p 0.533863mV 238018.438p 0.533863mV 238031.879p 0.551564mV 238045.778p 0.569279mV 238066.537p 0.604668mV 238078.881p 0.569858mV 238094.314p 0.587942mV 238098.781p 0.605667mV 239005.454p 0.56644mV 239025.235p 0.49616mV 239031.274p 0.513691mV 239053.638p 0.443164mV 240000.563p 0.551078mV 240024.839p 0.586171mV 240045.617p 0.568786mV 240058.297p 0.568976mV 240065.164p 0.534088mV 240085.248p 0.569653mV 240093.666p 0.552224mV 240098.735p 0.534814mV 240111.082p 0.552792mV 240125.827p 0.535722mV 240141.364p 0.553834mV 240145.361p 0.571576mV 241022.195p 0.546708mV 241043.509p 0.546674mV 241053.98p 0.581761mV 241087.178p 0.564468mV 241098.035p 0.564635mV 241103.975p 0.58228mV 241113.291p 0.617593mV 242013.852p 0.582397mV 242024.22p 0.582389mV 242028.068p 0.564855mV 242041.051p 0.547455mV 242049.819p 0.565086mV 242079.662p 0.565701mV 242122.489p 0.479779mV 242134.156p 0.515249mV 242153.966p 0.516096mV 243008.931p 0.56549mV 243015.564p 0.56557mV 243037.988p 0.6009mV 243068.117p 0.601656mV 244002.884p 0.552094mV 244007.241p 0.569595mV 244031.819p 0.622145mV 244057.431p 0.569971mV 244098.178p 0.536068mV 244122.823p 0.589412mV 245052.24p 0.515219mV 245063.501p 0.514991mV 245066.288p 0.532403mV 245070.117p 0.514706mV 245082.528p 0.51436mV 246056.037p 0.498188mV 246061.167p 0.515563mV 247021.769p 0.548725mV 247067.24p 0.530377mV 247074.321p 0.512696mV 247089.479p 0.494674mV 248014.565p 0.587283mV 248047.988p 0.605387mV 248059.918p 0.57061mV 248074.682p 0.588738mV 249018.922p 0.528664mV 249040.991p 0.475567mV 250046.001p 0.567337mV 250062.874p 0.584865mV 250091.86p 0.585056mV 250119.416p 0.567991mV 250128.892p 0.568257mV 250207.488p 0.501083mV 250208.78p 0.501083mV 250231.627p 0.484522mV 250271.923p 0.486157mV 251014.888p 0.550422mV 251017.271p 0.568048mV 251020.001p 0.585674mV 251026.577p 0.568194mV 251036.246p 0.533286mV 251043.257p 0.515842mV 251062.546p 0.481098mV 251119.676p 0.498897mV 251139.993p 0.428435mV 251142.586p 0.410781mV 252003.84p 0.553367mV 252024.164p 0.518367mV 252043.297p 0.5535mV 252068.748p 0.535848mV 252086.687p 0.500488mV 252087.714p 0.500488mV 253016.285p 0.4946mV 253061.773p 0.582095mV 253067.286p 0.599639mV 253091.092p 0.617437mV 253100.64p 0.582664mV 253101.475p 0.582664mV 253109.893p 0.600388mV 254005.47p 0.528143mV 254023.258p 0.545683mV 254033.069p 0.545684mV 254038.181p 0.528117mV 254042.433p 0.545673mV 254045.822p 0.563222mV 254070.383p 0.510536mV 254111.822p 0.474906mV 254112.584p 0.474906mV 254118.449p 0.492282mV 255006.684p 0.531204mV 255006.924p 0.531204mV 255023.429p 0.513567mV 255025.237p 0.531088mV 255028.344p 0.531088mV 255066.361p 0.530273mV 256048.637p 0.494799mV 256073.058p 0.582084mV 256077.44p 0.564417mV 256107.866p 0.528682mV 256114.406p 0.546116mV 256126.625p 0.563227mV 256176.988p 0.702431mV 256193.663p 0.75525mV 257003.118p 0.551889mV 257030.245p 0.586811mV 258004.975p 0.551798mV 258018.042p 0.534108mV 258019.246p 0.534108mV 258041.864p 0.516096mV 258065.931p 0.532753mV 258075.262p 0.49729mV 258079.323p 0.49729mV 259017.117p 0.529847mV 259108.839p 0.530276mV 259108.988p 0.530276mV 259152.175p 0.547915mV 259161.861p 0.583141mV 259194.275p 0.618907mV 260000.58p 0.553916mV 260012.017p 0.589092mV 260031.957p 0.659567mV 260042.802p 0.659828mV 261068.904p 0.534538mV 262008.782p 0.568941mV 262036.278p 0.53396mV 262058.695p 0.53416mV 262088.713p 0.499105mV 262100.163p 0.481299mV 262117.214p 0.428239mV 263027.812p 0.528789mV 263053.255p 0.546401mV 263055.909p 0.528859mV 263068.438p 0.528888mV 263087.793p 0.564019mV 263116.029p 0.599355mV 263116.844p 0.599355mV 263117.347p 0.599355mV 263135.457p 0.635056mV 263136.824p 0.635056mV 263138.826p 0.635056mV 264008.651p 0.531513mV 264019.819p 0.531399mV 264020.085p 0.513778mV 264024.285p 0.513778mV 264058.835p 0.56573mV 264078.326p 0.635479mV 264091.332p 0.582647mV 264093.326p 0.582647mV 264095.111p 0.600187mV 264112.103p 0.582604mV 264151.421p 0.582798mV 264178.469p 0.565421mV 264192.798p 0.583153mV 264220.564p 0.653914mV 264225.867p 0.67159mV 264231.856p 0.68927mV 265037.105p 0.497748mV 265039.973p 0.497748mV 265085.021p 0.53169mV 265086.148p 0.53169mV 266016.975p 0.601249mV 267018.783p 0.495493mV 267033.736p 0.477911mV 267035.341p 0.495428mV 267050.102p 0.512706mV 267056.726p 0.495027mV 267077.507p 0.459294mV 268028.239p 0.527874mV 268048.337p 0.562753mV 268060.829p 0.580128mV 268077.348p 0.562418mV 268077.516p 0.562418mV 268080.664p 0.544823mV 268103.304p 0.509523mV 268113.89p 0.544472mV 268114.7p 0.544472mV 268144.796p 0.614028mV 268156.544p 0.596266mV 268173.269p 0.57856mV 268211.932p 0.507692mV 269014.18p 0.587233mV 269018.848p 0.56968mV 269019.375p 0.56968mV 269030.219p 0.552206mV 269051.842p 0.552297mV 269054.128p 0.552297mV 269070.126p 0.587468mV 269075.305p 0.605049mV 269085.995p 0.60514mV 270013.984p 0.512964mV 271011.342p 0.51478mV 271022.732p 0.549784mV 272002.577p 0.547451mV 272037.072p 0.565144mV 272037.079p 0.565144mV 272049.461p 0.530088mV 272075.23p 0.600599mV 272088.224p 0.600836mV 272088.566p 0.600836mV 272126.085p 0.53234mV 272126.843p 0.53234mV 272144.159p 0.515558mV 273061.787p 0.616437mV 273068.327p 0.598919mV 273076.48p 0.599079mV 273100.037p 0.617308mV 274015.641p 0.496335mV 275028.27p 0.498017mV 275039.373p 0.497895mV 275045.797p 0.532764mV 275051.431p 0.55016mV 275078.861p 0.56691mV 275089.325p 0.566585mV 276008.867p 0.571332mV 276033.262p 0.553558mV 276034.606p 0.553558mV 276035.875p 0.535957mV 276039.714p 0.535957mV 276045.331p 0.500743mV 276055.243p 0.50059mV 276069.054p 0.465245mV 277005.387p 0.569785mV 277046.422p 0.569898mV 277064.113p 0.587658mV 277071.341p 0.587852mV 277082.321p 0.588098mV 277098.074p 0.606114mV 278000.054p 0.545753mV 278015.236p 0.493045mV 279006.732p 0.531318mV 279045.799p 0.60159mV 279050.93p 0.619214mV 280038.326p 0.564657mV 280054.158p 0.512308mV 280060.783p 0.547607mV 280062.381p 0.547607mV 280083.099p 0.477726mV 280089.054p 0.460227mV 280094.332p 0.442701mV 280105.54p 0.460186mV 280114.269p 0.442544mV 281006.399p 0.570576mV 281009.511p 0.570576mV 281010.403p 0.588111mV 281013.344p 0.588111mV 281022.729p 0.55297mV 281030.627p 0.588103mV 281032.034p 0.588103mV 281034.838p 0.588103mV 281068.592p 0.570852mV 281078.027p 0.570977mV 281087.34p 0.606238mV 281150.092p 0.520598mV 281204.353p 0.522117mV 281209.43p 0.504806mV 281223.997p 0.487996mV 282020.159p 0.586271mV 282028.58p 0.568802mV 282046.994p 0.569247mV 282047.536p 0.569247mV 282060.237p 0.622264mV 282072.796p 0.622594mV 283029.064p 0.530425mV 283039.998p 0.530333mV 283052.839p 0.477446mV 284051.219p 0.479664mV 284080.46p 0.443832mV 285002.569p 0.548496mV 285033.062p 0.548173mV 285070.415p 0.547386mV 285070.739p 0.547386mV 286013.945p 0.589048mV 286014.576p 0.589048mV 286015.149p 0.571435mV 286034.087p 0.553765mV 286065.792p 0.571145mV 286070.119p 0.588728mV 286087.591p 0.641526mV 286096.923p 0.641709mV 287013.987p 0.586mV 287035.732p 0.533491mV 287044.348p 0.55111mV 287076.294p 0.604364mV 287081.981p 0.622046mV 288035.338p 0.532481mV 288058.231p 0.497576mV 289017.364p 0.566162mV 289033.785p 0.548679mV 289037.91p 0.531168mV 289059.312p 0.531363mV 289069.745p 0.531474mV 289087.111p 0.531603mV 289147.264p 0.566813mV 289169.309p 0.531878mV 289182.098p 0.549661mV 289190.639p 0.549826mV 289210.407p 0.550255mV 290017.327p 0.566594mV 290027.132p 0.566632mV 290045.871p 0.601968mV 290071.841p 0.585213mV 291025.023p 0.603983mV 291044.339p 0.621595mV 291055.35p 0.569204mV 291087.718p 0.605252mV 292008.99p 0.570508mV 292045.376p 0.605987mV 292056.018p 0.641346mV 293016.532p 0.498945mV 293024.29p 0.481381mV 293026.599p 0.498918mV 293058.249p 0.463118mV 294007.841p 0.53094mV 294036.907p 0.460271mV 294041.007p 0.442598mV 294043.271p 0.442598mV 295007.12p 0.565849mV 295014.492p 0.548274mV 295015.307p 0.56583mV 295025.701p 0.530707mV 295030.29p 0.51315mV 295037.255p 0.495586mV 296005.918p 0.567331mV 296011.384p 0.549832mV 296014.37p 0.549832mV 296081.983p 0.586588mV 296082.513p 0.586588mV 296085.249p 0.569291mV 297009.443p 0.52984mV 297034.754p 0.476733mV 298013.552p 0.587947mV 298055.669p 0.570399mV 298058.658p 0.570399mV 298081.747p 0.588094mV 298111.611p 0.588571mV 298117.664p 0.571132mV 298143.788p 0.554324mV 298186.373p 0.503454mV 298254.557p 0.418039mV 298281.679p 0.382885mV 299014.12p 0.587021mV 299014.804p 0.587021mV 299022.744p 0.551943mV 299034.55p 0.552017mV 299051.895p 0.587277mV 299084.829p 0.622939mV 299086.893p 0.640629mV 300005.761p 0.532232mV 300013.086p 0.549795mV 300025.329p 0.49709mV 300029.1p 0.49709mV 300042.684p 0.514512mV 300043.632p 0.514512mV 300071.608p 0.548846mV 301013.024p 0.583967mV 301050.293p 0.478264mV 301054.962p 0.478264mV 302009.452p 0.529355mV 302015.389p 0.494197mV 302039.61p 0.529076mV 303001.561p 0.553253mV 303009.879p 0.535743mV 303011.781p 0.518232mV 303012.372p 0.518232mV 303076.651p 0.570998mV 303144.076p 0.624731mV 304037.663p 0.459476mV 305021.215p 0.580789mV 305031.134p 0.580918mV 305041.141p 0.616203mV 305062.723p 0.581743mV 306006.968p 0.567844mV 306019.066p 0.567915mV 306021.574p 0.550413mV 306029.674p 0.532921mV 306055.564p 0.498034mV 306085.457p 0.4977mV 306089.025p 0.4977mV 306110.558p 0.584789mV 306114.059p 0.584789mV 306125.845p 0.637073mV 306145.757p 0.636971mV 306148.77p 0.636971mV 306150.805p 0.619481mV 306152.667p 0.619481mV 306172.491p 0.620024mV 307003.252p 0.549428mV 307035.233p 0.532163mV 307048.712p 0.532275mV 307049.496p 0.532275mV 307075.863p 0.602837mV 307079.347p 0.602837mV 307083.982p 0.58536mV 307093.332p 0.585593mV 307112.945p 0.58625mV 308034.529p 0.617966mV 308052.158p 0.653491mV 309048.786p 0.533408mV 309102.772p 0.516682mV 309112.361p 0.516859mV 309140.671p 0.482021mV 309158.927p 0.499494mV 310014.394p 0.551388mV 310031.696p 0.621576mV 310058.921p 0.604332mV 310071.497p 0.587194mV 311033.884p 0.447351mV 312022.33p 0.514702mV 312024.918p 0.514702mV 312050.432p 0.549168mV 312058.078p 0.56654mV 312062.26p 0.548831mV 312063.297p 0.548831mV 312072.22p 0.58356mV 312074.217p 0.58356mV 312087.235p 0.600595mV 312105.709p 0.670262mV 312106.533p 0.670262mV 312126.192p 0.670166mV 312137.924p 0.670309mV 312141.452p 0.687978mV 312144.571p 0.687978mV 313046.088p 0.568995mV 313064.457p 0.551616mV 313073.575p 0.551771mV 313083.589p 0.551914mV 313089.033p 0.534438mV 313092.462p 0.516965mV 313130.473p 0.517203mV 313136.217p 0.534706mV 313139.171p 0.534706mV 313164.587p 0.551878mV 313173.221p 0.551704mV 313175.041p 0.569182mV 314009.282p 0.528602mV 314013.746p 0.511001mV 314023.933p 0.546002mV 314025.157p 0.528368mV 314029.206p 0.528368mV 314060.042p 0.50991mV 314064.237p 0.50991mV 315002.479p 0.550725mV 315030.046p 0.586291mV 315040.385p 0.55153mV 315042.605p 0.55153mV 315047.808p 0.53418mV 315069.741p 0.499837mV 315069.784p 0.499837mV 315105.854p 0.430651mV 316034.885p 0.583167mV 316042.683p 0.548045mV 316044.372p 0.548045mV 316067.64p 0.600776mV 316068.679p 0.600776mV 317011.394p 0.511528mV 317034.992p 0.546623mV 317054.439p 0.476342mV 318001.803p 0.546229mV 318012.191p 0.51107mV 318031.022p 0.440624mV 319017.165p 0.534169mV 319041.331p 0.551417mV 319072.074p 0.621312mV 319076.799p 0.638856mV 319080.457p 0.656424mV 319082.493p 0.656424mV 320015.304p 0.566878mV 320016.077p 0.566878mV 320017.296p 0.566878mV 320018.774p 0.566878mV 320028.298p 0.566853mV 320030.32p 0.584421mV 320034.416p 0.584421mV 320069.959p 0.672713mV 321017.268p 0.566529mV 321055.177p 0.46131mV 321073.671p 0.47857mV 321082.118p 0.443172mV 322000.593p 0.547864mV 322033.263p 0.477253mV 322054.928p 0.511722mV 323026.1p 0.531234mV 323030.209p 0.513635mV 323041.911p 0.478412mV 324014.25p 0.552575mV 324017.149p 0.570105mV 324038.444p 0.570031mV 324063.404p 0.51729mV 324096.63p 0.569219mV 324144.776p 0.515157mV 325003.545p 0.546939mV 325019.733p 0.529225mV 325068.188p 0.563578mV 325096.563p 0.563206mV 325103.331p 0.545563mV 325147.166p 0.632228mV 325170.42p 0.614279mV 325180.542p 0.57908mV 325206.363p 0.526148mV 325213.352p 0.508483mV 325214.354p 0.508483mV 326022.01p 0.554021mV 326026.223p 0.536438mV 326034.169p 0.553974mV 326074.938p 0.518483mV 327024.503p 0.480229mV 327024.555p 0.480229mV 327058.766p 0.567805mV 327075.728p 0.602741mV 327084.582p 0.620311mV 327098.179p 0.638036mV 328026.253p 0.569357mV 328067.594p 0.604406mV 329005.309p 0.571876mV 329042.963p 0.554698mV 329061.125p 0.590064mV 329075.648p 0.537685mV 329104.541p 0.485557mV 329105.909p 0.503189mV 329106.879p 0.503189mV 330011.574p 0.518317mV 330047.912p 0.500373mV 330054.197p 0.517821mV 330057.85p 0.535236mV 330124.601p 0.585486mV 330142.38p 0.65486mV 330157.224p 0.671984mV 330161.564p 0.689439mV 330167.976p 0.706924mV 330182.438p 0.689351mV 330184.827p 0.689351mV 331000.505p 0.546075mV 331008.786p 0.528535mV 331016.268p 0.528572mV 331059.463p 0.458069mV 331071.818p 0.510211mV 332048.23p 0.529317mV 332087.908p 0.564223mV 332088.481p 0.564223mV 332090.558p 0.546629mV 332100.554p 0.546579mV 332115.612p 0.528934mV 332124.18p 0.511351mV 332125.544p 0.493762mV 332131.666p 0.47616mV 332136.997p 0.493656mV 332162.537p 0.475425mV 333016.926p 0.60638mV 333033.146p 0.624064mV 333034.247p 0.624064mV 333052.328p 0.659615mV 334018.707p 0.534475mV 334034.121p 0.551922mV 334036.444p 0.569445mV 334049.839p 0.569372mV 334059.622p 0.569333mV 334063.948p 0.586888mV 334082.164p 0.586967mV 334085.185p 0.604571mV 334100.178p 0.622342mV 334112.254p 0.657661mV 335055.053p 0.458244mV 336022.618p 0.516019mV 336026.688p 0.498395mV 337001.174p 0.551209mV 337001.713p 0.551209mV 337020.505p 0.551336mV 337065.517p 0.498928mV 337072.795p 0.516463mV 337083.41p 0.551478mV 337094.507p 0.551355mV 337109.907p 0.568725mV 337145.966p 0.4983mV 337177.336p 0.532947mV 337214.573p 0.549557mV 338008.902p 0.571502mV 338021.73p 0.553913mV 338022.999p 0.553913mV 338034.609p 0.518815mV 338049.805p 0.53634mV 338088.925p 0.535918mV 338096.199p 0.570886mV 338100.199p 0.588362mV 338103.523p 0.588362mV 338125.493p 0.500231mV 338151.91p 0.5171mV 339010.78p 0.585359mV 339038.193p 0.603207mV 339039.755p 0.603207mV 339072.261p 0.586608mV 339082.514p 0.552003mV 340000.533p 0.549402mV 340008.661p 0.566962mV 340022.542p 0.549419mV 340027.824p 0.53186mV 341023.384p 0.587237mV 341030.232p 0.587212mV 341044.805p 0.622382mV 341070.291p 0.622991mV 341070.48p 0.622991mV 342023.367p 0.58615mV 342031.379p 0.621467mV 342032.955p 0.621467mV 343029.68p 0.494252mV 343040.453p 0.511608mV 343087.695p 0.598402mV 343088.418p 0.598402mV 343093.853p 0.580762mV 343110.594p 0.510261mV 343129.063p 0.49239mV 344020.429p 0.546183mV 344045.464p 0.528465mV 344052.593p 0.545978mV 344073.505p 0.615997mV 344086.237p 0.598429mV 344112.821p 0.651484mV 344112.897p 0.651484mV 345001.581p 0.55252mV 345024.86p 0.517668mV 346017.803p 0.567736mV 346051.929p 0.620396mV 346069.207p 0.568029mV 346080.278p 0.586017mV 346091.564p 0.551343mV 347014.771p 0.54892mV 347050.989p 0.549183mV 347053.744p 0.549183mV 347059.006p 0.566741mV 347082.062p 0.584447mV 347095.595p 0.602276mV 347101.948p 0.584874mV 347112.151p 0.620292mV 348000.709p 0.554185mV 348011.557p 0.589247mV 348019.116p 0.571663mV 348036.12p 0.571647mV 348056.299p 0.60689mV 348116.179p 0.608436mV 349010.785p 0.580829mV 349025.988p 0.633635mV 349038.36p 0.633831mV 349051.677p 0.581782mV 350001.146p 0.545854mV 350009.276p 0.528306mV 350021.347p 0.581013mV 350031.098p 0.545935mV 350082.539p 0.581728mV 350082.877p 0.581728mV 351000.757p 0.553791mV 351015.1p 0.571182mV 351032.549p 0.623696mV 352034.558p 0.551555mV 352038.676p 0.569163mV 352049.246p 0.569273mV 352076.978p 0.5698mV 352112.728p 0.51823mV 352162.617p 0.448486mV 352177.667p 0.430622mV 352186.687p 0.465298mV 353023.416p 0.585165mV 353057.58p 0.568545mV 353106.735p 0.535297mV 353120.868p 0.518291mV 353121.467p 0.518291mV 353169.068p 0.467568mV 354017.313p 0.571511mV 354026.987p 0.536532mV 354042.236p 0.554304mV 354061.154p 0.484403mV 354072.658p 0.519605mV 355140.666p 0.583826mV 355167.763p 0.495414mV 356002.956p 0.55141mV 356013.588p 0.551477mV 356059.918p 0.604474mV 356060.239p 0.586974mV 356080.01p 0.62251mV 357011.596p 0.551294mV 357017.588p 0.533784mV 357020.05p 0.516274mV 357023.599p 0.516274mV 357031.988p 0.516343mV 357032.031p 0.516343mV 357046.099p 0.533876mV 357046.387p 0.533876mV 357075.813p 0.42811mV 358018.341p 0.536133mV 358018.488p 0.536133mV 358036.715p 0.465877mV 359007.165p 0.533747mV 359009.177p 0.533747mV 359042.81p 0.516232mV 359078.081p 0.498093mV 359078.458p 0.498093mV 360004.023p 0.548953mV 360021.442p 0.584337mV 361000.209p 0.547959mV 361012.939p 0.512867mV 361013.82p 0.512867mV 361032.712p 0.477718mV 361043.984p 0.47761mV 361049.423p 0.495061mV 362001.215p 0.546776mV 362005.032p 0.564279mV 362022.79p 0.511446mV 362045.989p 0.493391mV 362049.344p 0.493391mV 363000.553p 0.547136mV 363005.578p 0.564662mV 363041.006p 0.582045mV 363101.257p 0.51217mV 363166.613p 0.599356mV 363169.815p 0.599356mV 363183.138p 0.616725mV 363184.952p 0.616725mV 363185.098p 0.634281mV 363195.403p 0.59923mV 363206.063p 0.634511mV 363223.637p 0.65246mV 364005.068p 0.564854mV 364007.108p 0.564854mV 364020.353p 0.582301mV 364021.82p 0.582301mV 364038.093p 0.529648mV 364046.288p 0.494556mV 364062.822p 0.441801mV 365074.815p 0.510801mV 365079.718p 0.528291mV 365108.832p 0.527665mV 366017.858p 0.604675mV 366039.68p 0.569966mV 366073.185p 0.448118mV 366081.766p 0.483348mV 366092.555p 0.448245mV 367003.839p 0.549713mV 367015.591p 0.602483mV 367047.401p 0.567853mV 367065.387p 0.498167mV 367075.38p 0.498383mV 367085.451p 0.53364mV 367091.036p 0.516139mV 367108.297p 0.498727mV 367128.791p 0.463573mV 368020.002p 0.588897mV 368021.549p 0.588897mV 368023.744p 0.588897mV 368035.894p 0.53644mV 368037.124p 0.53644mV 368082.99p 0.554492mV 368116.583p 0.572518mV 368124.77p 0.555114mV 368128.097p 0.537731mV 368130.948p 0.520361mV 368132.749p 0.520361mV 368156.571p 0.608906mV 369018.13p 0.528241mV 369018.808p 0.528241mV 369023.481p 0.51065mV 369036.285p 0.457815mV 369039.192p 0.457815mV 370010.659p 0.588082mV 370035.088p 0.570837mV 370036.908p 0.570837mV 370071.338p 0.483718mV 371000.003p 0.552207mV 371007.378p 0.569816mV 371020.429p 0.552427mV 371030.212p 0.587656mV 371046.418p 0.570341mV 371054.862p 0.587992mV 372017.956p 0.528413mV 372029.128p 0.528555mV 372039.434p 0.528664mV 372046.18p 0.528743mV 372102.342p 0.652368mV 373060.586p 0.510428mV 373066.46p 0.492791mV 373075.877p 0.492582mV 373082.865p 0.474906mV 374032.338p 0.518797mV 374086.368p 0.639436mV 374123.861p 0.655971mV 374124.64p 0.655971mV 374127.192p 0.673446mV 374127.388p 0.673446mV 374147.991p 0.67338mV 374149.368p 0.67338mV 374165.501p 0.708856mV 374168.465p 0.708856mV 374172.573p 0.691471mV 375015.927p 0.565757mV 375027.928p 0.565713mV 375034.372p 0.548148mV 375050.001p 0.583302mV 375058.285p 0.60089mV 375081.88p 0.653978mV 376002.618p 0.545523mV 376088.832p 0.527159mV 376098.714p 0.49179mV 377026.442p 0.568488mV 377056.615p 0.569161mV 377075.06p 0.499671mV 378063.24p 0.548193mV 378063.878p 0.548193mV 378073.022p 0.513417mV 378077.862p 0.531116mV 378097.817p 0.496619mV 378110.601p 0.5145mV 378136.381p 0.49743mV 378150.242p 0.480208mV 378150.743p 0.480208mV 378151.348p 0.480208mV 378169.088p 0.462959mV 379010.398p 0.583725mV 379030.407p 0.61884mV 379036.28p 0.601316mV 379107.443p 0.533033mV 379113.619p 0.550716mV 379118.028p 0.53331mV 379122.663p 0.551006mV 379133.758p 0.586406mV 380001.109p 0.547355mV 380018.743p 0.529623mV 380026.201p 0.564597mV 380052.185p 0.581876mV 380081.478p 0.546689mV 380099.744p 0.564219mV 380109.459p 0.599293mV 380110.953p 0.58172mV 380120.936p 0.581738mV 380129.223p 0.599329mV 380140.83p 0.617049mV 380146.077p 0.599575mV 380147.071p 0.599575mV 380166.469p 0.565003mV 380234.141p 0.478488mV 380247.84p 0.530923mV 380300.919p 0.582723mV 380327.623p 0.565066mV 380363.16p 0.617883mV 380365.176p 0.600424mV 381004.631p 0.54625mV 381058.6p 0.565008mV 382041.95p 0.479158mV 383036.96p 0.500731mV 383063.181p 0.447821mV 384000.306p 0.549629mV 384059.375p 0.426311mV 385027.871p 0.606565mV 385037.22p 0.641795mV 385048.315p 0.67709mV 385052.575p 0.694751mV 386005.906p 0.533444mV 386020.178p 0.551094mV 386028.006p 0.56869mV 386034.564p 0.551167mV 386035.049p 0.568772mV 386070.58p 0.481403mV 386092.018p 0.516531mV 386120.785p 0.551318mV 386173.463p 0.445173mV 387073.293p 0.476367mV 388012.826p 0.545994mV 388017.725p 0.528429mV 388026.385p 0.528417mV 388026.515p 0.528417mV 388086.067p 0.527414mV 388117.953p 0.561386mV 388118.632p 0.561386mV 388119.231p 0.561386mV 388120.811p 0.578753mV 389046.193p 0.564067mV 389049.553p 0.564067mV 389071.432p 0.582545mV 390004.712p 0.547999mV 390016.052p 0.565537mV 390030.397p 0.547945mV 390084.491p 0.618795mV 391004.388p 0.546544mV 391020.412p 0.511326mV 391033.99p 0.51124mV 391035.814p 0.493622mV 391050.614p 0.510895mV 391055.138p 0.528302mV 391079.668p 0.492526mV 392010.962p 0.584128mV 392011.871p 0.584128mV 392024.12p 0.584147mV 392033.955p 0.549122mV 393005.521p 0.569845mV 393038.054p 0.569754mV 393091.304p 0.658482mV 394004.822p 0.546305mV 394016.921p 0.56403mV 394017.672p 0.56403mV 394021.414p 0.581641mV 394026.255p 0.564143mV 394032.885p 0.546665mV 394052.985p 0.547053mV 394070.745p 0.582639mV 394101.65p 0.513734mV 394103.987p 0.513734mV 395018.437p 0.605093mV 395032.293p 0.587751mV 395039.717p 0.605416mV 396009.773p 0.532098mV 396029.05p 0.53193mV 396071.37p 0.478292mV 398018.881p 0.501043mV 398055.286p 0.570789mV 398060.416p 0.553163mV 398060.468p 0.553163mV 398087.509p 0.50013mV 398094.849p 0.517581mV 398104.791p 0.517305mV 398111.108p 0.551995mV 398111.549p 0.551995mV 398141.734p 0.550626mV 399003.521p 0.547317mV 399054.143p 0.582805mV 399058.172p 0.600468mV 399066.239p 0.600737mV 399070.933p 0.618436mV 400015.254p 0.533516mV 400027.799p 0.568457mV 400031.443p 0.58592mV 400033.924p 0.58592mV 400048.503p 0.568131mV 400056.611p 0.603093mV 400057.865p 0.603093mV 400069.446p 0.567866mV 400071.429p 0.585386mV 400128.145p 0.603339mV 401013.688p 0.548323mV 401028.666p 0.530866mV 401052.981p 0.618859mV 401059.385p 0.601374mV 401068.027p 0.56651mV 401080.096p 0.549444mV 401090.875p 0.514702mV 401103.969p 0.515037mV 401116.698p 0.533023mV 401141.85p 0.516169mV 401147.45p 0.53386mV 402008.446p 0.569849mV 402033.461p 0.552193mV 402037.295p 0.534634mV 402046.244p 0.534625mV 402056.789p 0.499473mV 402065.66p 0.534497mV 402084.224p 0.586904mV 402092.62p 0.551629mV 402134.084p 0.585918mV 402138.163p 0.56825mV 402140.355p 0.585689mV 402142.112p 0.585689mV 402144.922p 0.585689mV 402165.925p 0.567564mV 402170.865p 0.549905mV 402198.402p 0.49655mV 403031.373p 0.584331mV 403035.828p 0.601892mV 403040.541p 0.584344mV 403072.678p 0.549526mV 403092.836p 0.479458mV 403103.607p 0.514566mV 403130.39p 0.549317mV 403165.312p 0.531252mV 403165.718p 0.531252mV 403170.271p 0.513585mV 403189.254p 0.530702mV 403194.521p 0.548075mV 404012.645p 0.514531mV 404020.734p 0.514389mV 404052.192p 0.513592mV 405048.473p 0.60274mV 405091.387p 0.62084mV 406016.411p 0.533094mV 406033.037p 0.515309mV 406035.321p 0.497659mV 406109.048p 0.635983mV 406119.416p 0.600728mV 406122.904p 0.58312mV 406143.915p 0.653205mV 406144.679p 0.653205mV 406154.764p 0.653216mV 406167.478p 0.600727mV 406186.903p 0.566019mV 406189.727p 0.566019mV 406218.578p 0.601738mV 406232.593p 0.654816mV 406237.457p 0.637464mV 407006.978p 0.531017mV 407085.367p 0.530313mV 407102.66p 0.512238mV 407110.837p 0.511814mV 408015.744p 0.533834mV 408020.718p 0.551417mV 408020.928p 0.551417mV 408032.116p 0.55145mV 408061.553p 0.516342mV 408067.546p 0.533881mV 408067.671p 0.533881mV 408084.126p 0.55132mV 408087.525p 0.56883mV 408117.998p 0.568593mV 408123.126p 0.551mV 408125.403p 0.568534mV 408130.248p 0.586065mV 408133.968p 0.586065mV 408181.827p 0.621699mV 408185.603p 0.639385mV 409012.478p 0.519115mV 410062.096p 0.6165mV 410075.134p 0.669548mV 410078.38p 0.669548mV 410079.395p 0.669548mV 412015.481p 0.529541mV 412027.938p 0.529621mV 412033.127p 0.54722mV 412033.181p 0.54722mV 412044.329p 0.582412mV 412072.646p 0.582859mV 412092.182p 0.618481mV 412094.645p 0.618481mV 413036.494p 0.501908mV 413044.917p 0.519543mV 413184.307p 0.486487mV 413189.841p 0.504035mV 413196.078p 0.468861mV 413213.036p 0.486249mV 413215.51p 0.468603mV 414074.753p 0.586688mV 414079.675p 0.6042mV 414090.957p 0.621693mV 414118.959p 0.604371mV 414147.25p 0.570002mV 415028.303p 0.636981mV 415033.631p 0.654601mV 415041.536p 0.689891mV 415043.547p 0.689891mV 416001.228p 0.553674mV 416032.541p 0.48301mV 416059.599p 0.569845mV 416065.984p 0.569409mV 417014.086p 0.546299mV 417044.219p 0.475643mV 417048.223p 0.493079mV 418001.917p 0.54756mV 418002.313p 0.54756mV 418020.393p 0.547796mV 418048.991p 0.565721mV 418068.394p 0.566111mV 418075.047p 0.566358mV 418093.837p 0.584354mV 419055.443p 0.45975mV 420000.482p 0.551284mV 420010.712p 0.551232mV 420025.032p 0.533611mV 420049.921p 0.5686mV 420055.487p 0.568524mV 420060.131p 0.586063mV 420066.517p 0.568487mV 420095.967p 0.603729mV 420107.16p 0.603858mV 421065.897p 0.5272mV 421081.208p 0.544174mV 421104.287p 0.578318mV 422045.19p 0.59895mV 422065.142p 0.634565mV 423055.138p 0.568201mV 423070.311p 0.515962mV 423089.798p 0.463713mV 423098.457p 0.49899mV 424038.431p 0.465477mV 425035.527p 0.571241mV 425038.333p 0.571241mV 425060.779p 0.4841mV 425074.82p 0.484257mV 425104.365p 0.554531mV 426040.663p 0.588287mV 426057.491p 0.570485mV 426069.301p 0.53526mV 427001.842p 0.551789mV 427048.506p 0.498894mV 427056.208p 0.498637mV 427069.543p 0.49828mV 427069.905p 0.49828mV 428003.768p 0.547057mV 428009.64p 0.564627mV 428017.924p 0.564653mV 428029.763p 0.564723mV 428040.241p 0.547299mV 428056.667p 0.494741mV 429016.124p 0.536645mV 429042.555p 0.554235mV 429042.618p 0.554235mV 429043.267p 0.554235mV 429047.15p 0.571799mV 429048.831p 0.571799mV 429069.824p 0.642124mV 429089.344p 0.642574mV 430007.11p 0.53126mV 430020.035p 0.478506mV 430043.301p 0.443028mV 431003.018p 0.548558mV 431030.406p 0.548621mV 431053.942p 0.583665mV 431055.558p 0.601247mV 431098.525p 0.602151mV 432000.136p 0.546876mV 432001.562p 0.546876mV 432010.601p 0.546781mV 432018.304p 0.529167mV 432022.613p 0.511552mV 432024.643p 0.511552mV 432035.956p 0.528875mV 432070.957p 0.475271mV 433020.208p 0.5527mV 433051.334p 0.588468mV 434004.724p 0.54851mV 434015.509p 0.601299mV 434023.257p 0.618913mV 435007.427p 0.56398mV 435023.622p 0.581671mV 435067.31p 0.565406mV 436016.166p 0.570139mV 436112.327p 0.413185mV 436112.491p 0.413185mV 436121.434p 0.448059mV 436126.998p 0.430356mV 436128.745p 0.430356mV 437007.453p 0.535874mV 437016.147p 0.570938mV 437024.495p 0.588464mV 437029.059p 0.605997mV 437030.803p 0.623544mV 437036.959p 0.605988mV 437054.576p 0.623709mV 437069.177p 0.606523mV 438001.607p 0.55153mV 438005.156p 0.569147mV 438010.428p 0.551648mV 438013.378p 0.551648mV 438054.134p 0.587217mV 438067.228p 0.569866mV 438070.898p 0.552416mV 438082.4p 0.587752mV 438097.036p 0.605729mV 439035.146p 0.534964mV 439091.925p 0.552138mV 439095.593p 0.534503mV 439150.524p 0.621335mV 439159.772p 0.638867mV 439168.859p 0.674001mV 439174.14p 0.691607mV 440017.155p 0.530087mV 440020.905p 0.547686mV 440039.276p 0.600477mV 440079.56p 0.566344mV 440094.286p 0.549455mV 440095.979p 0.567209mV 441001.802p 0.550617mV 441008.205p 0.533106mV 441034.879p 0.515671mV 442015.284p 0.52829mV 442016.189p 0.52829mV 442017.806p 0.52829mV 442021.446p 0.510718mV 443019.384p 0.566901mV 443033.228p 0.549173mV 443041.671p 0.584151mV 443044.791p 0.584151mV 443059.657p 0.601542mV 444030.305p 0.549114mV 444055.404p 0.461541mV 444093.691p 0.548888mV 444096.987p 0.531229mV 444138.692p 0.635867mV 444143.46p 0.61829mV 444162.02p 0.618523mV 444170.588p 0.61883mV 444179.867p 0.601485mV 445006.48p 0.566509mV 445013.306p 0.548928mV 445021.545p 0.584023mV 445025.589p 0.601577mV 445037.725p 0.601614mV 445051.954p 0.584256mV 445063.119p 0.619596mV 446006.306p 0.563383mV 446015.687p 0.59851mV 446018.353p 0.59851mV 446056.258p 0.599249mV 446059.985p 0.599249mV 447032.48p 0.482066mV 447054.345p 0.551476mV 448002.269p 0.554358mV 448018.646p 0.607051mV 448029.256p 0.607121mV 448045.524p 0.642577mV 448045.844p 0.642577mV 448048.208p 0.642577mV 449025.534p 0.536447mV 449044.415p 0.588921mV 449149.817p 0.607945mV 450042.489p 0.443831mV 451017.337p 0.563756mV 451028.574p 0.528692mV 451047.375p 0.599054mV 451050.913p 0.616663mV 451061.57p 0.65193mV 451063.213p 0.65193mV 451063.678p 0.65193mV 452014.468p 0.549648mV 452018.36p 0.567255mV 452024.14p 0.549744mV 452071.941p 0.514961mV 452103.803p 0.479659mV 452125.943p 0.461497mV 452128.079p 0.461497mV 453006.226p 0.534221mV 453012.084p 0.551728mV 453124.967p 0.551546mV 453149.882p 0.604159mV 453152.884p 0.621722mV 454024.696p 0.623862mV 455022.019p 0.547563mV 455036.313p 0.530196mV 455059.824p 0.600672mV 455060.088p 0.618309mV 455077.016p 0.601152mV 456003.524p 0.553312mV 456043.728p 0.623687mV 456057.553p 0.641555mV 456060.053p 0.659244mV 456060.393p 0.659244mV 457000.394p 0.545862mV 457002.027p 0.545862mV 457002.447p 0.545862mV 457036.572p 0.598883mV 457054.183p 0.651923mV 458032.039p 0.550185mV 458032.128p 0.550185mV 458038.736p 0.532567mV 458041.933p 0.514947mV 458054.991p 0.51479mV 458062.449p 0.479456mV 459027.387p 0.599858mV 459038.444p 0.600006mV 459044.074p 0.617669mV 459044.102p 0.617669mV 460015.646p 0.501239mV 460043.485p 0.483524mV 461008.948p 0.53069mV 461011.914p 0.548202mV 461014.909p 0.548202mV 461032.49p 0.547984mV 461045.169p 0.495107mV 461065.39p 0.494584mV 462012.624p 0.546778mV 462015.067p 0.529245mV 462016.811p 0.529245mV 462020.347p 0.546831mV 462022.91p 0.546831mV 462074.883p 0.652952mV 463013.631p 0.583936mV 463015.128p 0.60149mV 463017.257p 0.60149mV 463058.791p 0.637241mV 464020.835p 0.546984mV 464025.044p 0.564594mV 464045.81p 0.599972mV 464046.231p 0.599972mV 465012.231p 0.581663mV 466037.209p 0.605386mV 466040.054p 0.623048mV 466047.977p 0.640721mV 467033.138p 0.580989mV 467038.235p 0.563461mV 467059.149p 0.598846mV 468002.962p 0.55398mV 468011.118p 0.553941mV 468012.251p 0.553941mV 468026.887p 0.606541mV 468030.291p 0.624093mV 469017.581p 0.493573mV 469038.801p 0.528585mV 469040.411p 0.510955mV 469042.117p 0.510955mV 470010.493p 0.514867mV 470071.421p 0.584623mV 470078.406p 0.60217mV 470081.57p 0.584607mV 470129.77p 0.603022mV 471068.298p 0.606338mV 471074.128p 0.589031mV 472052.698p 0.477025mV 473012.445p 0.514937mV 473021.098p 0.549936mV 473042.209p 0.514508mV 473053.887p 0.51431mV 474017.345p 0.564226mV 474033.201p 0.616962mV 474037.294p 0.63457mV 474047.706p 0.634745mV 475004.939p 0.550868mV 475036.518p 0.497927mV 475039.244p 0.497927mV 475066.173p 0.497336mV 475075.642p 0.497036mV 476006.013p 0.564303mV 476007.463p 0.564303mV 476028.295p 0.529112mV 476033.826p 0.511528mV 476048.333p 0.528955mV 476056.786p 0.563947mV 476079.256p 0.528553mV 476108.855p 0.527927mV 476110.705p 0.510245mV 478003.012p 0.548308mV 478026.665p 0.530663mV 478050.525p 0.583148mV 478051.419p 0.583148mV 478094.081p 0.618421mV 479014.588p 0.546111mV 479027.332p 0.528762mV 479048.562p 0.564164mV 479058.974p 0.599426mV 480000.637p 0.550571mV 480009.546p 0.533033mV 480029.129p 0.56824mV 480042.635p 0.585916mV 480049.733p 0.568419mV 480075.854p 0.63931mV 481017.31p 0.53333mV 481043.209p 0.58571mV 481049.939p 0.603231mV 481080.029p 0.621133mV 482010.114p 0.513216mV 482051.743p 0.478175mV 482082.918p 0.477349mV 483007.71p 0.568139mV 483027.123p 0.532904mV 483028.706p 0.532904mV 483030.666p 0.515294mV 484000.202p 0.553379mV 484013.358p 0.5533mV 484035.268p 0.535502mV 484080.726p 0.552223mV 484081.105p 0.552223mV 484100.717p 0.551763mV 484118.564p 0.568888mV 484136.885p 0.568163mV 484141.122p 0.585495mV 484176.444p 0.566394mV 485001.221p 0.550019mV 485004.383p 0.550019mV 485006.329p 0.567545mV 485035.428p 0.567366mV 485064.971p 0.54975mV 485065.608p 0.532165mV 485086.677p 0.532039mV 485131.646p 0.619447mV 485136.874p 0.636999mV 485146.339p 0.637056mV 485164.364p 0.619845mV 486012.783p 0.551029mV 486016.563p 0.568638mV 486026.673p 0.603863mV 486030.605p 0.586377mV 486031.082p 0.586377mV 486047.04p 0.604269mV 487028.013p 0.495569mV 487050.952p 0.512488mV 487059.908p 0.494759mV 488003.82p 0.546102mV 488005.11p 0.528548mV 488025.975p 0.563654mV 488076.352p 0.564143mV 488091.426p 0.617202mV 488098.505p 0.6349mV 489000.555p 0.546779mV 489043.982p 0.546787mV 489094.36p 0.546619mV 489095.876p 0.564168mV 489111.332p 0.546574mV 489111.417p 0.546574mV 489147.966p 0.528712mV 489163.463p 0.546059mV 490015.63p 0.601133mV 490063.103p 0.548536mV 490063.613p 0.548536mV 490088.085p 0.496069mV 491009.318p 0.563333mV 491013.981p 0.580883mV 491038.339p 0.598608mV 491040.255p 0.616248mV 491058.462p 0.599097mV 492014.893p 0.586966mV 492023.838p 0.62211mV 492045.121p 0.604996mV 493009.924p 0.532824mV 493017.739p 0.497691mV 493027.818p 0.497619mV 494026.019p 0.56464mV 494044.51p 0.546971mV 494045.342p 0.529383mV 494051.025p 0.511794mV 494077.486p 0.42366mV 495011.358p 0.582547mV 495109.502p 0.531492mV 495130.619p 0.619602mV 496017.988p 0.564571mV 496021.887p 0.582081mV 496023.522p 0.582081mV 496057.878p 0.634782mV 497017.988p 0.565905mV 497041.971p 0.548567mV 497110.218p 0.515333mV 497117.277p 0.533059mV 497175.643p 0.429894mV 497192.125p 0.447728mV 497218.393p 0.465493mV 497219.41p 0.465493mV 497226.257p 0.465472mV 497232.824p 0.483004mV 497251.153p 0.447711mV 497269.944p 0.46498mV 497282.708p 0.44703mV 498009.869p 0.56623mV 498020.286p 0.583976mV 498032.832p 0.584156mV 498067.812p 0.497304mV 498128.343p 0.568905mV 499003.08p 0.550084mV 499017.542p 0.602644mV 499028.752p 0.637743mV 499038.27p 0.637821mV 499041.839p 0.655465mV 499047.176p 0.638033mV 499057.157p 0.603335mV 500014.542p 0.515497mV 500056.606p 0.46198mV 501001.89p 0.552434mV 501028.999p 0.604855mV 501061.994p 0.622735mV 501066.619p 0.640425mV 501079.348p 0.64078mV 502034.543p 0.549554mV 502050.82p 0.549388mV 502052.587p 0.549388mV 502053.886p 0.549388mV 502096.24p 0.531347mV 502111.242p 0.548502mV 502124.743p 0.548193mV 502156.945p 0.564434mV 502170.673p 0.546249mV 503005.669p 0.565464mV 503009.061p 0.565464mV 504000.43p 0.550777mV 504021.844p 0.550668mV 504030.394p 0.550613mV 504051.451p 0.550465mV 504054.06p 0.550465mV 504063.245p 0.585518mV 504066.047p 0.603048mV 504070.821p 0.585469mV 504074.907p 0.585469mV 504080.504p 0.620602mV 504099.221p 0.63831mV 505007.351p 0.56801mV 505008.307p 0.56801mV 505015.962p 0.603131mV 505020.46p 0.62071mV 505053.159p 0.62142mV 506053.636p 0.588782mV 506057.263p 0.571315mV 506066.954p 0.571534mV 506094.953p 0.589815mV 507013.112p 0.517588mV 507018.864p 0.535101mV 507078.332p 0.674993mV 507088.605p 0.675161mV 508010.428p 0.51428mV 508035.783p 0.461562mV 508047.832p 0.461362mV 509058.88p 0.463584mV 509067.417p 0.463457mV 509082.379p 0.445492mV 509082.502p 0.445492mV 510008.077p 0.532766mV 510015.727p 0.567986mV 510028.616p 0.568088mV 510041.384p 0.515604mV 510041.454p 0.515604mV 510044.436p 0.515604mV 510076.126p 0.533294mV 510089.475p 0.533234mV 510091.984p 0.55075mV 510100.027p 0.550657mV 510117.553p 0.603198mV 510129.531p 0.568057mV 510143.149p 0.550568mV 510164.685p 0.515513mV 510174.584p 0.515497mV 510204.11p 0.550434mV 510209.855p 0.567976mV 510224.98p 0.585515mV 510231.781p 0.620705mV 510237.042p 0.603208mV 510243.797p 0.585748mV 511003.871p 0.553913mV 511005.446p 0.571518mV 511016.224p 0.5365mV 511057.462p 0.501525mV 511074.834p 0.483789mV 511083.999p 0.483535mV 511088.774p 0.465831mV 512000.551p 0.547859mV 512009.417p 0.565384mV 512033.017p 0.582868mV 512051.35p 0.618077mV 512089.062p 0.566285mV 512093.073p 0.548943mV 512098.78p 0.531621mV 512099.485p 0.531621mV 512165.66p 0.464158mV 512172.231p 0.481832mV 512250.706p 0.482829mV 512251.227p 0.482829mV 512253.004p 0.482829mV 513026.067p 0.535745mV 513037.208p 0.535627mV 513069.419p 0.499869mV 513073.011p 0.517199mV 514002.841p 0.548085mV 514007.784p 0.565639mV 514008.052p 0.565639mV 514008.743p 0.565639mV 514038.698p 0.600956mV 514054.823p 0.583863mV 515001.256p 0.546626mV 515008.807p 0.5291mV 515012.692p 0.511574mV 515029.521p 0.494045mV 515043.656p 0.511422mV 515063.565p 0.510869mV 516017.032p 0.569103mV 516019.971p 0.569103mV 516061.354p 0.587636mV 516079.35p 0.535531mV 516116.008p 0.502197mV 516155.804p 0.468912mV 516159.423p 0.468912mV 516170.327p 0.522075mV 517005.97p 0.567724mV 517006.942p 0.567724mV 517012.438p 0.550157mV 517019.286p 0.532598mV 517061.484p 0.479318mV 517064.425p 0.479318mV 517068.493p 0.496662mV 519017.036p 0.571448mV 519039.423p 0.606521mV 519074.676p 0.554193mV 520020.29p 0.549503mV 520034.454p 0.549618mV 520064.863p 0.549985mV 521022.962p 0.550402mV 521027.567p 0.567989mV 521041.073p 0.585656mV 521058.123p 0.603421mV 521064.945p 0.621068mV 522006.397p 0.571379mV 522019.692p 0.60643mV 522025.23p 0.606423mV 523070.027p 0.588066mV 524003.253p 0.552737mV 524003.603p 0.552737mV 524024.064p 0.482329mV 524032.707p 0.447056mV 525004.404p 0.550148mV 525025.835p 0.497399mV 526004.969p 0.548617mV 526010.807p 0.513489mV 526046.584p 0.56598mV 526053.034p 0.548383mV 526091.47p 0.548379mV 526119.184p 0.601338mV 526129.91p 0.601576mV 526137.832p 0.636975mV 527012.419p 0.517593mV 527054.42p 0.481942mV 527054.735p 0.481942mV 528036.384p 0.534975mV 528043.102p 0.517384mV 528058.431p 0.569904mV 528081.65p 0.552mV 528105.928p 0.569067mV 528115.157p 0.603982mV 528174.788p 0.621716mV 528178.354p 0.639403mV 528181.399p 0.622025mV 528189.012p 0.60469mV 529000.03p 0.547313mV 529000.587p 0.547313mV 529035.124p 0.494453mV 529051.954p 0.476663mV 529058.677p 0.458995mV 530034.153p 0.510274mV 530044.664p 0.474987mV 531004.392p 0.553481mV 531009.341p 0.57105mV 531019.588p 0.535953mV 531057.266p 0.500992mV 531070.379p 0.55365mV 531072.012p 0.55365mV 531089.113p 0.500878mV 531108.694p 0.500561mV 532018.116p 0.563634mV 532024.032p 0.581238mV 532025.679p 0.56373mV 532077.263p 0.495117mV 532098.312p 0.530939mV 532147.309p 0.462426mV 532162.901p 0.445097mV 533070.595p 0.616459mV 533093.14p 0.651831mV 534023.054p 0.511624mV 534055.586p 0.423666mV 535025.432p 0.565155mV 535026.458p 0.565155mV 535052.653p 0.547709mV 535067.404p 0.565374mV 535087.32p 0.495406mV 535138.314p 0.460137mV 535147.164p 0.424796mV 536014.289p 0.54865mV 536020.142p 0.548658mV 536031.798p 0.548678mV 536060.352p 0.54886mV 536099.885p 0.566798mV 537001.2p 0.547348mV 537014.994p 0.547306mV 537031.435p 0.547286mV 537036.95p 0.564865mV 537046.654p 0.564907mV 537062.54p 0.547487mV 537095.634p 0.670884mV 538019.407p 0.567391mV 538038.64p 0.602421mV 538060.904p 0.585014mV 538067.62p 0.602649mV 538070.435p 0.620294mV 538080.377p 0.65562mV 539050.279p 0.58759mV 539069.128p 0.605497mV 539080.977p 0.588479mV 540008.731p 0.563121mV 540039.257p 0.52836mV 540061.193p 0.546024mV 540061.925p 0.546024mV 540062.507p 0.546024mV 540063.21p 0.546024mV 540065.578p 0.528483mV 540090.243p 0.546162mV 540105.009p 0.528684mV 540142.479p 0.581726mV 540152.035p 0.58198mV 540152.493p 0.58198mV 540158.846p 0.599671mV 541007.38p 0.570013mV 541025.213p 0.570229mV 541026.735p 0.570229mV 541032.241p 0.552722mV 541034.097p 0.552722mV 541048.971p 0.570472mV 541052.205p 0.588115mV 541053.966p 0.588115mV 541055.054p 0.570657mV 541082.224p 0.553795mV 541092.126p 0.554161mV 541100.736p 0.589604mV 542004.083p 0.553312mV 542020.97p 0.553127mV 542023.598p 0.553127mV 542060.571p 0.552811mV 542080.703p 0.482337mV 543019.486p 0.529802mV 543039.351p 0.529937mV 543074.902p 0.512394mV 543076.193p 0.494781mV 543079.846p 0.494781mV 543127.649p 0.598628mV 543129.091p 0.598628mV 543166.111p 0.667686mV 543177.277p 0.667599mV 543177.852p 0.667599mV 543193.686p 0.650181mV 543200.152p 0.650447mV 543209.716p 0.668146mV 544010.863p 0.5494mV 544016.189p 0.567015mV 544062.543p 0.549949mV 544080.947p 0.550261mV 544129.604p 0.603965mV 544133.793p 0.586615mV 545000.46p 0.549574mV 545012.409p 0.549583mV 545028.449p 0.567196mV 545040.02p 0.54973mV 545054.28p 0.549822mV 545058.323p 0.532305mV 545066.843p 0.567509mV 545106.24p 0.603152mV 545112.384p 0.58575mV 545116.778p 0.603458mV 545127.961p 0.568817mV 546050.745p 0.476752mV 548027.096p 0.605126mV 548030.121p 0.587545mV 548069.367p 0.500035mV 548085.021p 0.53522mV 548115.07p 0.53495mV 548142.04p 0.481684mV 549029.4p 0.528925mV 549040.9p 0.546361mV 549045.861p 0.563853mV 549049.13p 0.563853mV 549061.15p 0.581223mV 549083.612p 0.581158mV 549109.998p 0.669129mV 550000.302p 0.553825mV 550006.134p 0.571424mV 550051.461p 0.44866mV 550052.034p 0.44866mV 551019.359p 0.528776mV 551068.122p 0.422754mV 552004.657p 0.54824mV 552018.905p 0.53069mV 552019.192p 0.53069mV 552039.03p 0.495545mV 553005.746p 0.535524mV 553055.271p 0.570855mV 553090.561p 0.659067mV 553093.828p 0.659067mV 554019.296p 0.605423mV 554022.048p 0.622968mV 554041.208p 0.658273mV 554045.043p 0.640867mV 555009.453p 0.5314mV 555030.795p 0.478379mV 556001.958p 0.552047mV 556006.772p 0.534507mV 556022.149p 0.552108mV 556042.117p 0.517024mV 556063.246p 0.481742mV 556066.076p 0.464084mV 556075.895p 0.4638mV 557028.342p 0.533124mV 557053.962p 0.515539mV 558042.822p 0.518739mV 558047.619p 0.536233mV 559007.037p 0.565981mV 559022.059p 0.548362mV 559067.025p 0.565707mV 559070.877p 0.583241mV 559092.181p 0.618364mV 560031.286p 0.514045mV 560038.389p 0.496473mV 561002.224p 0.553063mV 561007.884p 0.535505mV 561049.347p 0.500121mV 561071.179p 0.481858mV 562013.723p 0.547921mV 562039.89p 0.495478mV 562085.611p 0.459902mV 563027.315p 0.536869mV 563029.221p 0.536869mV 563045.478p 0.571963mV 563059.765p 0.571938mV 563075.43p 0.607129mV 563105.162p 0.64283mV 563109.329p 0.64283mV 564026.144p 0.532587mV 564053.274p 0.479766mV 564079.103p 0.496699mV 564080.927p 0.478979mV 565030.933p 0.589603mV 565054.982p 0.625173mV 566000.084p 0.545974mV 566000.906p 0.545974mV 566053.603p 0.475583mV 567000.093p 0.546042mV 567004.166p 0.546042mV 567078.936p 0.563244mV 567079.212p 0.563244mV 567082.186p 0.580869mV 567101.165p 0.546096mV 567111.201p 0.54629mV 567119.298p 0.528843mV 567124.479p 0.511397mV 567137.812p 0.52921mV 567150.226p 0.511824mV 567161.494p 0.511928mV 567174.106p 0.547129mV 567196.561p 0.600106mV 567198.233p 0.600106mV 568045.809p 0.498887mV 568069.815p 0.463248mV 569005.43p 0.53173mV 569031.932p 0.478882mV 569039.359p 0.496364mV 569048.247p 0.531224mV 569060.818p 0.5132mV 570016.019p 0.565109mV 570032.56p 0.617826mV 570054.907p 0.618128mV 570057.459p 0.635796mV 571019.315p 0.570214mV 571063.994p 0.623479mV 571064.178p 0.623479mV 571065.914p 0.606111mV 571068.363p 0.606111mV 572065.475p 0.634169mV 572066.523p 0.634169mV 572075.294p 0.63435mV 572087.302p 0.599619mV 573007.827p 0.531363mV 573041.784p 0.549067mV 573065.325p 0.63683mV 573069.416p 0.63683mV 574038.572p 0.568996mV 574064.976p 0.516626mV 574087.419p 0.534354mV 574097.439p 0.534361mV 574111.294p 0.481627mV 574114.307p 0.481627mV 574122.477p 0.481514mV 574147.892p 0.498386mV 575015.789p 0.571824mV 575016.763p 0.571824mV 575020.371p 0.589441mV 575025.42p 0.607063mV 575051.28p 0.660301mV 576002.05p 0.550267mV 576019.275p 0.532708mV 576020.994p 0.550251mV 576023.376p 0.550251mV 576038.76p 0.602869mV 576056.298p 0.567869mV 576092.51p 0.550919mV 576093.922p 0.550919mV 576158.932p 0.499353mV 576177.486p 0.534499mV 576201.749p 0.481813mV 576220.182p 0.481645mV 577021.537p 0.519156mV 577030.39p 0.519067mV 577061.348p 0.553514mV 577076.54p 0.570603mV 577083.416p 0.552901mV 577155.466p 0.567371mV 577158.522p 0.567371mV 578013.72p 0.546967mV 578038.213p 0.529158mV 578054.124p 0.511423mV 578084.791p 0.475522mV 579057.119p 0.496096mV 579061.38p 0.478526mV 579078.648p 0.4608mV 579081.357p 0.478224mV 579094.232p 0.477875mV 580027.897p 0.534733mV 580039.483p 0.534807mV 580056.233p 0.464643mV 580101.448p 0.551467mV 580126.935p 0.568474mV 580148.813p 0.533013mV 580161.002p 0.515057mV 580166.608p 0.532434mV 580185.25p 0.531585mV 581064.185p 0.510721mV 581093.012p 0.509891mV 581094.553p 0.509891mV 582038.736p 0.52955mV 582040.098p 0.546942mV 582040.601p 0.546942mV 583007.949p 0.568779mV 583012.187p 0.551274mV 583040.81p 0.481247mV 583042.865p 0.481247mV 584036.542p 0.564802mV 584041.653p 0.547173mV 584045.631p 0.564664mV 584060.645p 0.546908mV 584079.957p 0.529103mV 585002.344p 0.550897mV 585005.372p 0.568472mV 585017.304p 0.603627mV 585018.637p 0.603627mV 585050.263p 0.586698mV 586011.025p 0.550438mV 586018.528p 0.568054mV 586024.698p 0.58567mV 587034.073p 0.549814mV 587039.816p 0.56739mV 587057.45p 0.567486mV 587068.019p 0.56756mV 587078.915p 0.567682mV 587109.028p 0.56825mV 587112.379p 0.550842mV 587163.78p 0.552445mV 587179.545p 0.500546mV 587184.074p 0.518301mV 587188.564p 0.536054mV 588038.202p 0.599719mV 588047.534p 0.599911mV 588050.076p 0.617581mV 588064.305p 0.652947mV 589003.123p 0.549337mV 589016.325p 0.531904mV 589023.765p 0.549503mV 589052.46p 0.620091mV 589065.142p 0.568019mV 590002.526p 0.550051mV 590016.15p 0.567683mV 590057.448p 0.603703mV 591018.683p 0.534763mV 591057.545p 0.534807mV 591062.0p 0.552393mV 591067.469p 0.534852mV 591106.278p 0.570157mV 591112.702p 0.552633mV 591116.458p 0.53512mV 591126.591p 0.535215mV 591142.636p 0.588036mV 591156.103p 0.640929mV 591167.31p 0.641189mV 592001.276p 0.550196mV 592038.575p 0.638042mV 592052.82p 0.585666mV 592081.609p 0.586791mV 593003.065p 0.553457mV 593006.883p 0.535857mV 593047.113p 0.500199mV 593060.062p 0.482209mV 593061.246p 0.482209mV 594012.472p 0.547121mV 594023.851p 0.547018mV 594024.366p 0.547018mV 594032.209p 0.511777mV 594033.135p 0.511777mV 594055.979p 0.528776mV 594066.643p 0.493366mV 594070.02p 0.475655mV 595009.005p 0.56987mV 595073.781p 0.587309mV 595079.342p 0.569856mV 595084.753p 0.552421mV 595086.821p 0.570093mV 595097.37p 0.605439mV 595117.948p 0.606111mV 596026.903p 0.535679mV 596041.717p 0.517912mV 596041.795p 0.517912mV 597028.244p 0.497649mV 597038.467p 0.532828mV 597082.799p 0.550373mV 597087.352p 0.567905mV 597112.158p 0.585381mV 597123.75p 0.585389mV 597139.381p 0.568001mV 597142.721p 0.550546mV 597182.016p 0.5517mV 598013.498p 0.549786mV 598042.556p 0.549988mV 598044.748p 0.549988mV 598066.095p 0.462348mV 599033.568p 0.581699mV 599043.364p 0.546738mV 599056.861p 0.49436mV 599083.244p 0.512115mV 599093.744p 0.512064mV 599101.42p 0.476844mV 600011.806p 0.588837mV 600042.99p 0.589035mV 600069.762p 0.572148mV 600079.77p 0.537426mV 600081.596p 0.555148mV 600082.1p 0.555148mV 600102.61p 0.591009mV 601002.491p 0.550259mV 601003.049p 0.550259mV 601017.907p 0.532645mV 601044.144p 0.51498mV 601073.936p 0.54966mV 601082.042p 0.584594mV 601124.488p 0.61955mV 603040.558p 0.51346mV 604017.919p 0.569095mV 604030.25p 0.586836mV 604044.368p 0.622146mV 605011.803p 0.580882mV 605071.014p 0.51069mV 605109.749p 0.562886mV 605146.154p 0.668178mV 606021.2p 0.582755mV 606035.974p 0.530116mV 606043.713p 0.512581mV 606068.722p 0.530025mV 606111.284p 0.546466mV 606116.252p 0.563879mV 606128.223p 0.563595mV 606162.593p 0.54484mV 607009.258p 0.566227mV 607030.612p 0.654109mV 608011.328p 0.514133mV 608028.23p 0.531738mV 608035.079p 0.496588mV 608051.454p 0.47887mV 608099.716p 0.59991mV 608119.062p 0.564043mV 608135.905p 0.563226mV 609006.157p 0.565454mV 609019.586p 0.565479mV 609078.532p 0.636677mV 610012.317p 0.580839mV 610016.481p 0.563227mV 610022.039p 0.545626mV 610029.907p 0.563149mV 610051.907p 0.580591mV 611038.202p 0.603532mV 611042.684p 0.621143mV 611047.49p 0.638771mV 612027.496p 0.534992mV 612054.646p 0.482042mV 613032.982p 0.514426mV 614003.062p 0.551222mV 614032.814p 0.516265mV 615035.831p 0.53616mV 616021.733p 0.547199mV 616027.769p 0.564794mV 616081.198p 0.477634mV 616095.196p 0.460121mV 616111.646p 0.477456mV 616116.539p 0.494871mV 616130.619p 0.511884mV 616145.79p 0.563771mV 616153.347p 0.546017mV 616153.807p 0.546017mV 616158.306p 0.563297mV 617002.846p 0.551407mV 617009.233p 0.533813mV 617041.285p 0.551003mV 617047.877p 0.568511mV 617048.282p 0.568511mV 617095.887p 0.46226mV 618005.324p 0.530225mV 618088.05p 0.566337mV 618092.414p 0.548934mV 618113.523p 0.549649mV 618122.897p 0.585134mV 619005.64p 0.531353mV 619011.249p 0.513842mV 619029.075p 0.496357mV 619058.525p 0.460739mV 620000.663p 0.551404mV 620003.597p 0.551404mV 620014.999p 0.516242mV 620033.29p 0.516062mV 620039.378p 0.533531mV 620050.494p 0.515653mV 620060.928p 0.515394mV 621023.815p 0.550114mV 621071.432p 0.620352mV 622002.615p 0.548602mV 622007.741p 0.530984mV 622053.567p 0.618334mV 622057.669p 0.600774mV 622080.168p 0.618708mV 622090.022p 0.619051mV 622092.488p 0.619051mV 623016.22p 0.563473mV 623071.012p 0.511038mV 623107.594p 0.563227mV 623108.195p 0.563227mV 623116.365p 0.563097mV 623185.269p 0.59871mV 624000.401p 0.54828mV 624037.151p 0.530771mV 624044.063p 0.548325mV 624051.487p 0.5483mV 624079.531p 0.60098mV 624104.351p 0.583829mV 625037.046p 0.634138mV 625043.753p 0.616601mV 625056.532p 0.634405mV 625069.897p 0.634729mV 626000.099p 0.545724mV 626005.294p 0.528156mV 626009.171p 0.528156mV 626049.46p 0.633553mV 626052.752p 0.616062mV 626068.979p 0.669056mV 627007.002p 0.569829mV 627098.194p 0.570238mV 627107.394p 0.570497mV 627111.044p 0.553091mV 627145.899p 0.53666mV 627155.081p 0.536995mV 627163.366p 0.554703mV 628003.203p 0.54784mV 628005.312p 0.565435mV 628071.967p 0.477174mV 628075.268p 0.49452mV 629003.368p 0.546493mV 629028.679p 0.493598mV 629029.154p 0.493598mV 630003.932p 0.548624mV 630038.397p 0.636534mV 631015.42p 0.529171mV 631019.803p 0.529171mV 631030.548p 0.581724mV 631038.69p 0.599243mV 631046.983p 0.634331mV 631058.769p 0.634397mV 631070.165p 0.652244mV 631073.017p 0.652244mV 631078.901p 0.669935mV 632127.63p 0.53192mV 632172.941p 0.478377mV 633059.634p 0.498993mV 634022.211p 0.620189mV 634024.837p 0.620189mV 634027.878p 0.602689mV 634042.575p 0.585468mV 635006.244p 0.536057mV 635020.923p 0.518572mV 635035.212p 0.46588mV 635049.177p 0.500862mV 636000.141p 0.549836mV 636013.921p 0.514755mV 636039.624p 0.49704mV 636048.656p 0.496832mV 637045.752p 0.531375mV 637079.593p 0.565417mV 637112.212p 0.581446mV 637120.214p 0.580965mV 638003.52p 0.550995mV 638020.221p 0.515993mV 638066.391p 0.427726mV 639005.325p 0.532909mV 639017.535p 0.532983mV 639030.17p 0.585713mV 639047.612p 0.603398mV 639049.182p 0.603398mV 640042.201p 0.581699mV 641014.556p 0.58568mV 641019.882p 0.568129mV 641020.691p 0.585712mV 641023.495p 0.585712mV 641024.15p 0.585712mV 641030.087p 0.620903mV 641086.059p 0.53441mV 641089.239p 0.53441mV 642005.212p 0.531948mV 642031.972p 0.584456mV 642042.557p 0.619516mV 642049.187p 0.601952mV 642055.26p 0.566898mV 642066.762p 0.5319mV 642078.029p 0.496893mV 642083.255p 0.479367mV 642115.441p 0.531607mV 643011.597p 0.581859mV 643012.388p 0.581859mV 643028.079p 0.599601mV 644024.286p 0.549901mV 644052.108p 0.549732mV 644081.444p 0.549353mV 644085.735p 0.566859mV 644090.746p 0.549243mV 644112.765p 0.584139mV 644119.235p 0.60165mV 644120.807p 0.584051mV 644138.73p 0.566434mV 644152.865p 0.54884mV 644176.709p 0.531062mV 644197.419p 0.565751mV 644201.616p 0.548087mV 644201.824p 0.548087mV 644217.565p 0.600352mV 644224.73p 0.582671mV 644225.248p 0.564995mV 644234.245p 0.582416mV 644246.634p 0.59955mV 644249.234p 0.59955mV 644279.927p 0.563601mV 645013.671p 0.51617mV 645013.945p 0.51617mV 645018.458p 0.533699mV 645029.817p 0.533595mV 645053.784p 0.48044mV 646016.908p 0.530662mV 646021.779p 0.51313mV 646026.931p 0.530712mV 646034.607p 0.513158mV 646057.542p 0.460292mV 646068.746p 0.460061mV 647138.285p 0.60411mV 647141.059p 0.586794mV 648012.646p 0.51349mV 648028.41p 0.495868mV 648039.385p 0.46065mV 648054.008p 0.477859mV 649023.79p 0.583602mV 649044.003p 0.583561mV 649086.718p 0.531229mV 649088.069p 0.531229mV 649103.708p 0.513762mV 649149.544p 0.495753mV 649164.424p 0.51281mV 649182.717p 0.546986mV 649189.049p 0.564261mV 650020.325p 0.551246mV 650047.213p 0.568504mV 650070.734p 0.620845mV 650080.636p 0.655939mV 650081.375p 0.655939mV 650093.93p 0.65602mV 650094.57p 0.65602mV 650103.43p 0.656244mV 651019.022p 0.568957mV 651020.638p 0.586543mV 651060.448p 0.587415mV 652003.206p 0.548502mV 652015.229p 0.5659mV 652030.642p 0.583301mV 652065.868p 0.671368mV 653001.192p 0.546968mV 653008.688p 0.564529mV 653058.927p 0.458905mV 654020.805p 0.588828mV 654043.813p 0.624225mV 655008.498p 0.531673mV 655060.666p 0.584654mV 655062.938p 0.584654mV 655071.51p 0.584743mV 655080.23p 0.584886mV 655085.044p 0.602544mV 655092.398p 0.62021mV 655105.862p 0.603171mV 655106.699p 0.603171mV 656022.264p 0.582917mV 656052.944p 0.61876mV 657050.552p 0.551084mV 657054.364p 0.551084mV 657055.457p 0.533449mV 657081.711p 0.515394mV 658003.802p 0.550691mV 658022.58p 0.515602mV 658038.931p 0.533137mV 658052.845p 0.51546mV 659039.693p 0.599311mV 659056.872p 0.56466mV 659056.915p 0.56466mV 659069.718p 0.529887mV 659073.343p 0.512511mV 659076.618p 0.495131mV 659089.387p 0.495412mV 659090.195p 0.513086mV 660005.975p 0.566839mV 660011.605p 0.549307mV 660025.185p 0.531848mV 660064.829p 0.549236mV 660083.458p 0.619252mV 660116.062p 0.672194mV 660116.345p 0.672194mV 661009.675p 0.529518mV 661064.441p 0.581644mV 661064.649p 0.581644mV 661082.602p 0.651687mV 661086.675p 0.634138mV 661089.164p 0.634138mV 661093.778p 0.616627mV 662001.201p 0.547814mV 662014.148p 0.582982mV 662037.318p 0.530563mV 662046.682p 0.530694mV 662058.615p 0.530792mV 662077.003p 0.530945mV 662128.209p 0.460082mV 662132.162p 0.477443mV 663005.244p 0.570231mV 663049.996p 0.64109mV 664005.793p 0.528611mV 664029.104p 0.458131mV 664041.222p 0.440191mV 665006.314p 0.564278mV 665007.603p 0.564278mV 665028.082p 0.564456mV 665039.922p 0.564644mV 665041.072p 0.547194mV 665070.325p 0.477598mV 665081.547p 0.477682mV 665100.43p 0.51274mV 665141.88p 0.47705mV 665156.724p 0.529297mV 665189.444p 0.598335mV 665198.881p 0.598007mV 665200.037p 0.615401mV 665202.957p 0.615401mV 665246.333p 0.667821mV 665257.364p 0.703152mV 666007.438p 0.529153mV 666083.247p 0.4757mV 667006.107p 0.56362mV 667021.016p 0.616366mV 668006.63p 0.57197mV 668028.781p 0.571977mV 668039.739p 0.536911mV 668137.895p 0.570278mV 668144.288p 0.58759mV 668150.315p 0.552113mV 668172.343p 0.586222mV 668176.76p 0.603475mV 669015.435p 0.564767mV 669037.986p 0.599793mV 669048.293p 0.634926mV 669062.863p 0.617579mV 670027.625p 0.493974mV 670056.987p 0.528381mV 670063.575p 0.545705mV 670065.725p 0.563013mV 670074.137p 0.580312mV 671046.586p 0.564319mV 671108.767p 0.49522mV 671121.608p 0.442845mV 671124.557p 0.442845mV 671132.163p 0.478029mV 671140.41p 0.477996mV 671151.366p 0.477875mV 671180.104p 0.477064mV 672013.607p 0.551228mV 672032.495p 0.621459mV 672044.77p 0.656667mV 673035.145p 0.533227mV 673058.003p 0.497639mV 673075.127p 0.567013mV 673078.744p 0.567013mV 673088.671p 0.531515mV 674007.65p 0.569096mV 674016.743p 0.5341mV 674048.796p 0.464028mV 674062.43p 0.481376mV 674071.443p 0.446014mV 675001.932p 0.551677mV 675022.216p 0.551432mV 675042.877p 0.586345mV 675087.459p 0.639338mV 675089.653p 0.639338mV 675099.202p 0.639631mV 676049.54p 0.534982mV 676052.224p 0.552423mV 676061.43p 0.552173mV 676074.184p 0.586977mV 676087.567p 0.604116mV 676098.634p 0.568811mV 676103.615p 0.586276mV 676154.583p 0.550474mV 676189.673p 0.567041mV 676189.847p 0.567041mV 677002.317p 0.552814mV 677011.711p 0.517749mV 677041.668p 0.552687mV 677044.35p 0.552687mV 677088.131p 0.534061mV 678006.816p 0.565334mV 678017.402p 0.565352mV 678018.721p 0.565352mV 678024.888p 0.547802mV 678077.38p 0.566027mV 678082.977p 0.548652mV 678088.258p 0.566366mV 678095.662p 0.566735mV 678112.92p 0.514802mV 678129.573p 0.533009mV 678163.937p 0.482184mV 678168.917p 0.499945mV 679023.084p 0.545433mV 679036.264p 0.56282mV 679036.439p 0.56282mV 679042.416p 0.545205mV 679063.411p 0.544964mV 679070.594p 0.509687mV 679084.613p 0.474381mV 680023.797p 0.552609mV 680025.682p 0.53508mV 680028.469p 0.53508mV 680048.689p 0.57031mV 680075.841p 0.53566mV 680101.778p 0.553756mV 680147.179p 0.467457mV 680155.779p 0.432626mV 682016.728p 0.563781mV 682022.862p 0.546208mV 682025.904p 0.528642mV 682047.012p 0.56371mV 682048.481p 0.56371mV 682055.829p 0.528551mV 682066.399p 0.52851mV 682107.96p 0.52806mV 682118.85p 0.527871mV 682162.787p 0.50904mV 682163.29p 0.50904mV 683029.931p 0.602082mV 683040.089p 0.619859mV 684022.227p 0.588734mV 684023.927p 0.588734mV 684091.526p 0.589812mV 685032.598p 0.548023mV 685058.863p 0.565398mV 685073.54p 0.582913mV 685074.477p 0.582913mV 685085.268p 0.600486mV 685095.618p 0.600601mV 685127.385p 0.566166mV 685137.576p 0.531387mV 685165.706p 0.497205mV 685167.304p 0.497205mV 685174.14p 0.514888mV 685190.582p 0.51539mV 685245.209p 0.499049mV 685247.107p 0.499049mV 685280.698p 0.552315mV 685282.409p 0.552315mV 685287.567p 0.569963mV 686013.788p 0.51816mV 686018.327p 0.535723mV 686056.541p 0.535226mV 686066.472p 0.534917mV 686077.951p 0.499489mV 687058.039p 0.496771mV 687061.371p 0.514239mV 687070.034p 0.513999mV 687074.107p 0.513999mV 688003.738p 0.552951mV 688013.209p 0.517881mV 688021.827p 0.517899mV 688031.867p 0.517843mV 688041.157p 0.517743mV 688042.466p 0.517743mV 688078.088p 0.534326mV 689005.975p 0.53508mV 689011.898p 0.517496mV 689026.54p 0.499796mV 689040.897p 0.481945mV 689046.486p 0.499326mV 690005.127p 0.531058mV 690009.023p 0.531058mV 690012.603p 0.513551mV 690063.236p 0.548376mV 690068.985p 0.530755mV 690090.852p 0.547914mV 690171.039p 0.618006mV 691052.901p 0.652005mV 691054.372p 0.652005mV 692036.47p 0.600787mV 692060.12p 0.54912mV 692080.965p 0.515102mV 692091.17p 0.515588mV 693049.0p 0.424349mV 694005.658p 0.5363mV 694013.53p 0.518682mV 694020.585p 0.518533mV 694047.745p 0.46528mV 695000.859p 0.549847mV 695007.171p 0.567356mV 695018.784p 0.532143mV 695051.945p 0.549202mV 695057.432p 0.531554mV 695059.897p 0.531554mV 695082.2p 0.478325mV 696005.093p 0.535907mV 696012.255p 0.553488mV 696016.94p 0.535941mV 696053.109p 0.483281mV 696063.558p 0.483186mV 696075.832p 0.465329mV 696080.022p 0.447649mV 697019.199p 0.566902mV 697040.275p 0.584802mV 697041.154p 0.584802mV 697049.218p 0.602448mV 697065.615p 0.567912mV 697075.606p 0.603352mV 697083.82p 0.621075mV 698032.273p 0.512574mV 698057.364p 0.494453mV 698065.739p 0.494151mV 699017.966p 0.499991mV 700020.68p 0.515854mV 701017.961p 0.563096mV 701029.053p 0.56302mV 701035.016p 0.56298mV 701038.816p 0.56298mV 701064.855p 0.545312mV 701079.818p 0.562748mV 701086.962p 0.562666mV 701124.527p 0.509642mV 701143.796p 0.439033mV 702010.444p 0.516869mV 702012.554p 0.516869mV 702026.981p 0.534402mV 702055.375p 0.604432mV 702066.022p 0.604475mV 702069.756p 0.604475mV 702071.394p 0.622079mV 702081.563p 0.657338mV 702087.594p 0.639899mV 702091.262p 0.657587mV 703010.582p 0.55083mV 703032.78p 0.515952mV 703035.571p 0.533561mV 703046.575p 0.568748mV 703072.321p 0.551515mV 703109.423p 0.570066mV 703114.18p 0.587777mV 703114.648p 0.587777mV 704005.184p 0.567254mV 704041.466p 0.479857mV 705013.217p 0.554418mV 705018.165p 0.571992mV 705021.79p 0.589565mV 705030.57p 0.58962mV 705032.093p 0.58962mV 705078.991p 0.537503mV 705085.407p 0.502538mV 705086.036p 0.502538mV 705122.525p 0.555182mV 705136.604p 0.607688mV 705155.371p 0.607717mV 705169.851p 0.572745mV 705180.601p 0.555542mV 705211.594p 0.556277mV 705224.264p 0.521409mV 705238.857p 0.574436mV 706044.877p 0.550193mV 706054.283p 0.550285mV 706062.73p 0.58549mV 706068.606p 0.567984mV 706074.363p 0.550499mV 706076.831p 0.533027mV 706081.317p 0.55067mV 706111.913p 0.516154mV 706151.889p 0.587299mV 706161.394p 0.552613mV 707041.803p 0.581215mV 707043.14p 0.581215mV 707048.653p 0.598818mV 707067.564p 0.599173mV 707078.532p 0.564429mV 708002.759p 0.552401mV 708043.193p 0.587241mV 708047.267p 0.604814mV 708095.213p 0.535109mV 708146.666p 0.499329mV 708160.811p 0.516264mV 709004.48p 0.550702mV 709004.652p 0.550702mV 709027.093p 0.497818mV 709034.484p 0.515303mV 709035.638p 0.497653mV 709047.215p 0.497413mV 709049.795p 0.497413mV 709061.931p 0.514439mV 709066.755p 0.53174mV 710023.035p 0.51189mV 710029.257p 0.52948mV 710034.311p 0.511937mV 710034.471p 0.511937mV 710042.753p 0.51195mV 710070.896p 0.546897mV 710077.672p 0.564396mV 710127.373p 0.528965mV 710143.859p 0.581522mV 710154.684p 0.616581mV 710175.589p 0.599239mV 710182.584p 0.616893mV 710186.567p 0.599462mV 711008.793p 0.535012mV 711016.42p 0.534948mV 711025.546p 0.569955mV 711055.34p 0.640026mV 711062.364p 0.657621mV 711067.936p 0.675239mV 712012.32p 0.581033mV 712024.25p 0.581124mV 712049.278p 0.564069mV 712080.129p 0.477348mV 712100.219p 0.512731mV 712127.81p 0.495267mV 712171.399p 0.547334mV 712175.27p 0.564819mV 712178.553p 0.564819mV 712183.819p 0.547201mV 712207.985p 0.564647mV 712213.099p 0.547086mV 712243.158p 0.547425mV 712258.703p 0.530273mV 712258.795p 0.530273mV 712267.923p 0.565641mV 712270.397p 0.583331mV 712279.722p 0.601028mV 714022.619p 0.581201mV 714029.207p 0.56363mV 714034.507p 0.546076mV 714048.711p 0.563673mV 714066.535p 0.563743mV 714082.909p 0.616575mV 714089.449p 0.634211mV 714092.045p 0.651864mV 714103.366p 0.617092mV 715020.502p 0.547875mV 715020.975p 0.547875mV 715044.324p 0.477435mV 715057.469p 0.494654mV 716000.29p 0.553534mV 716030.929p 0.588794mV 717001.754p 0.554344mV 717031.766p 0.484155mV 717052.833p 0.518981mV 717056.165p 0.501294mV 718033.228p 0.621932mV 718043.839p 0.621971mV 718054.938p 0.622125mV 719009.612p 0.530395mV 719041.222p 0.58249mV 719093.367p 0.546384mV 720057.762p 0.459428mV 720078.485p 0.49419mV 720092.68p 0.511193mV 721002.308p 0.546941mV 721007.779p 0.529332mV 721018.697p 0.564339mV 721028.525p 0.529107mV 721033.98p 0.511492mV 722015.721p 0.568022mV 722038.937p 0.638341mV 722066.504p 0.569043mV 722068.458p 0.569043mV 722074.196p 0.586791mV 723032.039p 0.514945mV 724000.142p 0.549832mV 724002.332p 0.549832mV 724025.72p 0.532191mV 724051.073p 0.51421mV 725014.009p 0.550208mV 725017.529p 0.567807mV 725020.219p 0.585405mV 725038.171p 0.568042mV 725075.757p 0.533993mV 725084.556p 0.551669mV 725100.212p 0.552225mV 726018.963p 0.601999mV 727050.679p 0.510729mV 728001.403p 0.546514mV 728019.521p 0.529119mV 728051.651p 0.546873mV 728053.071p 0.546873mV 728055.998p 0.529328mV 728066.123p 0.529358mV 728096.958p 0.529185mV 728112.225p 0.546471mV 728117.024p 0.528811mV 728130.288p 0.546007mV 728175.82p 0.597597mV 728212.196p 0.614814mV 728214.328p 0.614814mV 728229.976p 0.63245mV 728244.757p 0.650237mV 728247.043p 0.632833mV 728259.716p 0.668251mV 729000.284p 0.547521mV 729021.383p 0.582699mV 729027.868p 0.565155mV 729029.636p 0.565155mV 729041.541p 0.582837mV 730000.284p 0.55186mV 730010.349p 0.516616mV 730054.714p 0.585579mV 730059.173p 0.6029mV 730125.65p 0.671384mV 730130.869p 0.688955mV 730160.948p 0.689608mV 731030.034p 0.549283mV 731040.079p 0.514199mV 731048.435p 0.496649mV 731069.078p 0.531612mV 732006.008p 0.570566mV 732009.114p 0.570566mV 732023.005p 0.588147mV 733005.918p 0.531345mV 733080.615p 0.512801mV 733088.112p 0.53013mV 734031.794p 0.550359mV 734044.491p 0.55011mV 734073.797p 0.514196mV 735024.677p 0.550438mV 735026.177p 0.567919mV 735055.225p 0.637762mV 735062.979p 0.655309mV 735073.168p 0.690486mV 735081.469p 0.690666mV 735082.23p 0.690666mV 736000.367p 0.550758mV 736017.344p 0.603612mV 736043.132p 0.656803mV 737022.671p 0.549085mV 737043.359p 0.478928mV 737055.669p 0.496381mV 737062.377p 0.51385mV 737064.769p 0.51385mV 737085.283p 0.495565mV 738017.155p 0.536613mV 738029.545p 0.501357mV 738048.878p 0.571082mV 738063.09p 0.588187mV 738084.339p 0.517433mV 739021.616p 0.547535mV 739028.116p 0.565045mV 739107.423p 0.598897mV 739122.1p 0.616231mV 739146.029p 0.63368mV 739165.221p 0.598878mV 739182.021p 0.616827mV 739200.233p 0.582523mV 740004.957p 0.553555mV 740017.321p 0.536034mV 740079.936p 0.570781mV 740080.445p 0.553161mV 740104.025p 0.517774mV 741024.317p 0.589801mV 741027.173p 0.607422mV 741041.683p 0.625264mV 741060.872p 0.590902mV 741062.796p 0.590902mV 742027.195p 0.570025mV 742027.236p 0.570025mV 742068.176p 0.605459mV 742076.308p 0.605753mV 743012.425p 0.581347mV 743035.929p 0.56408mV 743045.727p 0.529135mV 743056.13p 0.494207mV 743108.543p 0.494806mV 743161.168p 0.442315mV 744033.893p 0.585663mV 744036.01p 0.568154mV 744043.253p 0.585777mV 745110.811p 0.586603mV 745117.333p 0.604281mV 746007.314p 0.536098mV 746029.218p 0.571074mV 746036.611p 0.571039mV 746043.701p 0.588583mV 746047.11p 0.571011mV 746075.074p 0.571145mV 746085.933p 0.60638mV 746144.756p 0.590177mV 746146.374p 0.607893mV 746151.807p 0.590565mV 747003.979p 0.550137mV 747011.368p 0.515075mV 747020.587p 0.550224mV 747022.344p 0.550224mV 747023.729p 0.550224mV 747037.435p 0.567794mV 747043.278p 0.585379mV 747048.904p 0.567851mV 747076.806p 0.603459mV 747096.123p 0.56905mV 748004.765p 0.554079mV 748023.116p 0.589248mV 748030.311p 0.554176mV 748039.166p 0.571777mV 748069.634p 0.607386mV 749015.448p 0.605584mV 749021.678p 0.623206mV 750019.228p 0.606751mV 750025.208p 0.571722mV 750144.855p 0.554253mV 750152.942p 0.554133mV 750154.164p 0.554133mV 750175.556p 0.501059mV 751037.426p 0.532262mV 751048.697p 0.532112mV 751067.137p 0.566809mV 751109.608p 0.4956mV 752017.342p 0.533796mV 753016.516p 0.532612mV 753040.07p 0.585101mV 753064.053p 0.585022mV 753081.519p 0.620309mV 753108.72p 0.6385mV 754054.856p 0.545919mV 754066.78p 0.563556mV 754121.141p 0.546841mV 754153.384p 0.512525mV 754154.938p 0.512525mV 754156.768p 0.495121mV 754158.029p 0.495121mV 754173.091p 0.513037mV 754178.678p 0.49558mV 755016.363p 0.601526mV 755018.111p 0.601526mV 755021.599p 0.584002mV 755026.118p 0.601619mV 755069.616p 0.602739mV 756012.794p 0.551356mV 756065.355p 0.60482mV 757009.916p 0.56875mV 757018.308p 0.603931mV 757034.226p 0.621691mV 757045.639p 0.604544mV 757046.07p 0.604544mV 758010.545p 0.5524mV 758014.294p 0.5524mV 758017.665p 0.569919mV 758037.647p 0.604944mV 758040.788p 0.622517mV 758042.137p 0.622517mV 758067.543p 0.675577mV 758067.704p 0.675577mV 759011.982p 0.546759mV 759047.641p 0.529442mV 759082.406p 0.441496mV 760002.188p 0.547096mV 760005.196p 0.564714mV 760019.017p 0.56484mV 760049.093p 0.565367mV 760073.056p 0.513454mV 760078.782p 0.531143mV 760123.366p 0.514461mV 761041.014p 0.615958mV 762009.465p 0.536343mV 762013.117p 0.553904mV 762013.162p 0.553904mV 762024.147p 0.58901mV 762028.92p 0.571448mV 762050.994p 0.62433mV 762052.246p 0.62433mV 762056.368p 0.641992mV 762072.261p 0.624953mV 763013.554p 0.545952mV 763020.06p 0.545987mV 763025.668p 0.563557mV 763031.139p 0.581127mV 763038.403p 0.598704mV 763063.78p 0.546347mV 763085.697p 0.56448mV 763166.296p 0.460506mV 764028.225p 0.495068mV 764033.795p 0.477519mV 764045.757p 0.459857mV 764065.708p 0.529409mV 764066.12p 0.529409mV 764078.556p 0.564006mV 764093.792p 0.545789mV 765017.946p 0.500471mV 765056.592p 0.50011mV 766035.088p 0.532332mV 766078.306p 0.462158mV 767004.149p 0.547577mV 767029.425p 0.529896mV 767031.109p 0.51231mV 767035.728p 0.529836mV 767043.091p 0.547343mV 767043.861p 0.547343mV 767079.774p 0.529088mV 767084.2p 0.511392mV 768005.335p 0.564519mV 768019.547p 0.564607mV 768025.525p 0.529595mV 768044.796p 0.512201mV 768078.981p 0.565149mV 768088.247p 0.565291mV 768164.468p 0.444203mV 769095.304p 0.565026mV 769098.252p 0.565026mV 769103.22p 0.582625mV 769133.806p 0.618338mV 770008.184p 0.535206mV 770052.076p 0.482754mV 771033.586p 0.480208mV 771035.357p 0.497634mV 772045.625p 0.56327mV 772049.857p 0.56327mV 772051.548p 0.580898mV 772060.945p 0.581068mV 772062.34p 0.581068mV 772064.813p 0.581068mV 772069.595p 0.563635mV 773018.676p 0.571071mV 773036.22p 0.571078mV 773072.067p 0.518859mV 773083.952p 0.554108mV 773125.302p 0.572651mV 774008.259p 0.563395mV 774020.962p 0.51059mV 774023.252p 0.51059mV 774036.65p 0.527973mV 774052.695p 0.580361mV 774075.814p 0.632763mV 775005.053p 0.563602mV 775009.453p 0.563602mV 775028.448p 0.528508mV 775028.739p 0.528508mV 775033.376p 0.546075mV 775049.485p 0.528524mV 775066.838p 0.493394mV 775105.425p 0.562609mV 775114.984p 0.544882mV 775123.305p 0.544489mV 776001.559p 0.547801mV 776031.1p 0.547385mV 776035.838p 0.564871mV 776037.583p 0.564871mV 776063.836p 0.547013mV 776090.958p 0.511393mV 776112.37p 0.510731mV 776116.11p 0.49301mV 777015.28p 0.496522mV 777119.224p 0.706584mV 778033.836p 0.516777mV 778053.878p 0.551726mV 778064.348p 0.516515mV 778074.392p 0.516388mV 778085.989p 0.533604mV 778110.205p 0.515271mV 779008.822p 0.533334mV 779021.529p 0.515616mV 779022.847p 0.515616mV 779027.15p 0.497994mV 779038.578p 0.497815mV 779044.766p 0.480139mV 779048.745p 0.462453mV 780007.231p 0.570801mV 780009.371p 0.570801mV 781002.26p 0.547179mV 781010.391p 0.51194mV 781012.573p 0.51194mV 781050.006p 0.510854mV 782007.645p 0.531307mV 782058.188p 0.60197mV 782077.473p 0.567609mV 782084.027p 0.585345mV 783043.315p 0.585033mV 783055.482p 0.637625mV 783059.576p 0.637625mV 783093.125p 0.620693mV 784010.64p 0.585395mV 784030.53p 0.585691mV 784033.194p 0.585691mV 784059.978p 0.568793mV 785038.267p 0.600981mV 786029.437p 0.571211mV 786073.701p 0.482831mV 787004.984p 0.553039mV 787007.267p 0.535474mV 787022.203p 0.517869mV 787025.904p 0.50026mV 787035.737p 0.535221mV 787043.284p 0.552667mV 788010.693p 0.552705mV 788013.487p 0.552705mV 788027.007p 0.535149mV 788051.565p 0.517559mV 789001.004p 0.548578mV 789003.019p 0.548578mV 789037.99p 0.565753mV 789054.939p 0.583221mV 789056.383p 0.600782mV 789061.162p 0.618355mV 789082.219p 0.583494mV 789122.799p 0.549382mV 789135.191p 0.532143mV 789186.038p 0.427269mV 790016.316p 0.530816mV 790046.359p 0.566292mV 791029.001p 0.534218mV 791041.201p 0.55176mV 791055.719p 0.604405mV 792024.344p 0.58944mV 792026.441p 0.571863mV 792035.882p 0.536741mV 792044.996p 0.554304mV 792049.181p 0.571858mV 792057.072p 0.571846mV 792154.922p 0.591343mV 793027.623p 0.601585mV 793034.564p 0.584134mV 794041.633p 0.54577mV 794045.847p 0.528184mV 795017.81p 0.57006mV 795054.127p 0.623325mV 796058.801p 0.568922mV 796070.198p 0.586316mV 796090.783p 0.586228mV 796097.266p 0.568669mV 796105.823p 0.603812mV 796161.323p 0.516703mV 796178.36p 0.534454mV 796218.014p 0.569683mV 796232.835p 0.58726mV 796295.803p 0.499922mV 796305.001p 0.499976mV 796311.564p 0.517528mV 797023.412p 0.476299mV 797048.665p 0.563978mV 797057.688p 0.563883mV 797073.248p 0.581385mV 797096.909p 0.564009mV 797101.444p 0.581625mV 797108.33p 0.564131mV 797164.999p 0.512824mV 797166.937p 0.495407mV 797174.793p 0.477982mV 797175.442p 0.460541mV 797200.874p 0.408019mV 798006.49p 0.566058mV 798017.352p 0.601055mV 798053.994p 0.618631mV 798071.676p 0.584037mV 798084.518p 0.584428mV 799003.27p 0.550055mV 799011.238p 0.550059mV 799015.833p 0.532491mV 799018.571p 0.532491mV 799025.139p 0.532471mV 799041.726p 0.549926mV 799048.585p 0.567438mV 799100.11p 0.585376mV 800045.572p 0.565197mV 800078.736p 0.634854mV 800116.112p 0.599891mV 800137.842p 0.635463mV 800144.591p 0.65315mV 801008.426p 0.535089mV 801037.404p 0.534784mV 801057.705p 0.464168mV 802014.627p 0.55447mV 802022.574p 0.554538mV 802023.782p 0.554538mV 802034.474p 0.554598mV 802067.184p 0.572656mV 802083.595p 0.590629mV 802093.265p 0.626044mV 803014.987p 0.547158mV 803016.941p 0.56467mV 803022.433p 0.582183mV 803031.83p 0.617241mV 803058.882p 0.600006mV 804007.378p 0.529952mV 804078.346p 0.493743mV 805007.546p 0.533516mV 805013.587p 0.51596mV 805024.265p 0.480819mV 805050.022p 0.410095mV 806022.043p 0.547475mV 806033.84p 0.547526mV 806062.43p 0.477361mV 806062.557p 0.477361mV 806073.477p 0.477256mV 806076.238p 0.459605mV 807000.658p 0.549399mV 807013.518p 0.514343mV 807045.365p 0.496459mV 807053.096p 0.513837mV 808041.011p 0.550181mV 808045.544p 0.532634mV 809006.519p 0.536679mV 809070.629p 0.589951mV 809108.672p 0.538049mV 809125.818p 0.503531mV 809180.036p 0.522346mV 809208.028p 0.575769mV 810018.956p 0.56783mV 810021.287p 0.550278mV 810029.788p 0.532732mV 810040.165p 0.550323mV 811006.138p 0.569934mV 811055.968p 0.500492mV 811082.005p 0.447831mV 811082.057p 0.447831mV 812024.046p 0.552015mV 812052.79p 0.552275mV 812074.943p 0.517272mV 812091.439p 0.552369mV 812097.212p 0.534798mV 812104.441p 0.517231mV 813040.859p 0.58117mV 813053.363p 0.546169mV 813069.647p 0.493721mV 813082.406p 0.511401mV 813122.376p 0.616614mV 813154.186p 0.652206mV 814019.463p 0.567383mV 814022.391p 0.584979mV 814067.439p 0.603538mV 814074.479p 0.586197mV 815012.402p 0.552253mV 815030.671p 0.587595mV 815035.29p 0.60522mV 815061.383p 0.553207mV 815106.506p 0.572259mV 815109.776p 0.572259mV 815114.355p 0.554868mV 816047.93p 0.565226mV 816077.419p 0.635401mV 816087.873p 0.635522mV 817006.608p 0.569477mV 817022.819p 0.587242mV 817030.827p 0.552362mV 817056.992p 0.500312mV 817087.266p 0.500707mV 817106.798p 0.465716mV 817139.743p 0.535641mV 817145.573p 0.535455mV 817203.614p 0.551892mV 817221.99p 0.516375mV 817270.342p 0.549752mV 817281.668p 0.549341mV 818012.607p 0.581499mV 818030.905p 0.651739mV 818030.964p 0.651739mV 818033.689p 0.651739mV 818041.092p 0.686988mV 819059.358p 0.534913mV 820005.866p 0.52914mV 820006.154p 0.52914mV 820010.858p 0.54673mV 820016.394p 0.564313mV 820042.702p 0.617222mV 820046.469p 0.599764mV 820048.254p 0.599764mV 820049.187p 0.599764mV 820067.281p 0.530251mV 821010.58p 0.551976mV 822029.984p 0.49892mV 823007.586p 0.536548mV 823009.079p 0.536548mV 823014.444p 0.518988mV 823025.725p 0.501354mV 823031.285p 0.518837mV 823062.261p 0.517967mV 823066.504p 0.535266mV 824024.08p 0.548859mV 824052.184p 0.51331mV 824058.514p 0.530781mV 824081.998p 0.47748mV 825075.56p 0.570291mV 825095.952p 0.535501mV 825099.779p 0.535501mV 825122.048p 0.518409mV 825190.194p 0.517892mV 825224.54p 0.516539mV 826000.514p 0.547944mV 826069.951p 0.600139mV 826086.681p 0.635431mV 826094.403p 0.653072mV 827010.058p 0.550828mV 827039.364p 0.603441mV 827068.676p 0.568649mV 827104.417p 0.551969mV 827113.838p 0.587335mV 828025.293p 0.528065mV 828081.41p 0.580195mV 828113.697p 0.509828mV 828124.853p 0.509785mV 828150.216p 0.544402mV 828159.579p 0.561804mV 828185.219p 0.525776mV 828188.048p 0.525776mV 829021.042p 0.587757mV 829055.963p 0.570067mV 829073.992p 0.552456mV 829083.628p 0.517337mV 829107.912p 0.464423mV 829110.931p 0.446748mV 830029.179p 0.571978mV 830043.065p 0.554572mV 830092.64p 0.625552mV 831040.931p 0.658253mV 832010.443p 0.550549mV 832031.879p 0.515606mV 832090.223p 0.550342mV 832091.961p 0.550342mV 833013.132p 0.515694mV 833019.168p 0.533187mV 833019.638p 0.533187mV 833037.621p 0.46259mV 833040.819p 0.444915mV 834007.623p 0.563622mV 834017.87p 0.563645mV 834028.175p 0.528589mV 834069.744p 0.599207mV 835000.108p 0.5544mV 835023.91p 0.519159mV 835029.638p 0.536647mV 835033.749p 0.554117mV 835045.817p 0.536276mV 835060.557p 0.518401mV 836056.431p 0.641234mV 836060.008p 0.623739mV 836065.695p 0.64139mV 836070.185p 0.623963mV 836073.651p 0.623963mV 837040.538p 0.582173mV 838020.901p 0.551686mV 838027.728p 0.534102mV 838045.833p 0.56912mV 838052.37p 0.551553mV 838057.292p 0.533993mV 838076.2p 0.604223mV 838080.218p 0.621798mV 839010.069p 0.583349mV 839022.98p 0.618385mV 839046.145p 0.706362mV 840005.925p 0.529651mV 840013.691p 0.547178mV 840024.488p 0.547095mV 840061.178p 0.582106mV 840074.231p 0.61736mV 840085.866p 0.600174mV 840086.174p 0.600174mV 840095.742p 0.600556mV 841002.865p 0.550646mV 841010.082p 0.515486mV 841028.447p 0.497805mV 841045.052p 0.462237mV 842004.271p 0.550388mV 842019.64p 0.602908mV 842021.614p 0.585315mV 842030.92p 0.585303mV 842043.538p 0.620479mV 842055.682p 0.603154mV 842063.609p 0.585719mV 842068.006p 0.603403mV 842080.728p 0.621437mV 842088.887p 0.639153mV 843000.543p 0.552264mV 843001.45p 0.552264mV 843020.107p 0.516991mV 843023.581p 0.516991mV 843051.198p 0.551477mV 843061.119p 0.551149mV 843061.213p 0.551149mV 843090.373p 0.58499mV 843095.571p 0.60229mV 843105.459p 0.566806mV 844013.583p 0.517455mV 844020.645p 0.517453mV 844025.519p 0.499876mV 844039.619p 0.534913mV 844061.123p 0.51696mV 844068.453p 0.49931mV 845016.651p 0.53424mV 845061.95p 0.550834mV 845066.745p 0.568178mV 845086.295p 0.602444mV 845107.631p 0.531546mV 845111.053p 0.548865mV 846019.385p 0.529526mV 846019.418p 0.529526mV 846068.739p 0.565173mV 846069.331p 0.565173mV 846078.557p 0.565434mV 846082.381p 0.548027mV 846083.336p 0.548027mV 846089.295p 0.565722mV 846108.953p 0.531326mV 846109.304p 0.531326mV 846115.594p 0.496642mV 846150.677p 0.515261mV 846187.971p 0.463401mV 846188.449p 0.463401mV 846214.346p 0.44601mV 846238.045p 0.428205mV 846239.85p 0.428205mV 847000.691p 0.551029mV 847011.32p 0.551027mV 847013.585p 0.551027mV 848011.103p 0.55221mV 848018.035p 0.569806mV 848044.038p 0.622756mV 849017.127p 0.496161mV 849030.394p 0.478532mV 849047.637p 0.530939mV 849050.011p 0.513261mV 849052.879p 0.513261mV 849070.758p 0.51264mV 849078.566p 0.494922mV 850034.947p 0.482244mV 850059.604p 0.499231mV 851010.306p 0.547395mV 851024.103p 0.582381mV 851034.258p 0.547159mV 851116.956p 0.564912mV 851131.389p 0.582592mV 851152.134p 0.547744mV 852026.503p 0.566551mV 852048.422p 0.496315mV 852056.29p 0.496257mV 852066.958p 0.531236mV 852111.665p 0.582768mV 852125.647p 0.599938mV 852128.076p 0.599938mV 852138.702p 0.634831mV 852147.961p 0.634695mV 852162.4p 0.617127mV 852186.375p 0.63509mV 853038.848p 0.637797mV 853042.556p 0.655437mV 853043.506p 0.655437mV 853043.927p 0.655437mV 853044.691p 0.655437mV 853049.554p 0.638002mV 854005.878p 0.529643mV 854016.334p 0.494438mV 854020.059p 0.476822mV 854034.844p 0.476645mV 855012.176p 0.552652mV 855023.457p 0.55255mV 855024.282p 0.55255mV 855024.66p 0.55255mV 855080.187p 0.551323mV 855088.216p 0.568726mV 855128.846p 0.532192mV 856010.874p 0.517432mV 856011.916p 0.517432mV 856035.167p 0.535059mV 856077.135p 0.534996mV 856078.628p 0.534996mV 856088.924p 0.499829mV 856100.959p 0.517196mV 856123.078p 0.551713mV 856123.581p 0.551713mV 856139.504p 0.568674mV 856161.504p 0.585209mV 856165.833p 0.602579mV 856172.1p 0.619951mV 856198.121p 0.601693mV 856207.044p 0.566326mV 856208.524p 0.566326mV 856221.652p 0.618484mV 856232.688p 0.618146mV 856237.708p 0.635511mV 856244.614p 0.652878mV 856260.29p 0.652281mV 856275.439p 0.669439mV 856279.419p 0.669439mV 856290.072p 0.686772mV 856294.38p 0.686772mV 856320.133p 0.686956mV 856323.767p 0.686956mV 857017.891p 0.535023mV 857023.832p 0.517481mV 857034.785p 0.482369mV 858000.384p 0.553307mV 858013.22p 0.518183mV 858016.377p 0.535736mV 858026.343p 0.570804mV 858028.006p 0.570804mV 858035.001p 0.535632mV 858049.09p 0.535581mV 858066.245p 0.500282mV 858072.15p 0.517764mV 858118.563p 0.533916mV 859007.785p 0.529924mV 859015.288p 0.530044mV 859020.226p 0.512527mV 859030.576p 0.547708mV 859058.936p 0.530277mV 859108.072p 0.494811mV 859111.969p 0.477121mV 859116.257p 0.494496mV 860038.26p 0.564597mV 860061.948p 0.582271mV 860071.255p 0.617554mV 860079.92p 0.635213mV 860088.626p 0.635502mV 861014.387p 0.554278mV 861015.467p 0.571837mV 861084.826p 0.590134mV 861091.461p 0.555452mV 862019.454p 0.492901mV 862025.076p 0.457722mV 863001.981p 0.546144mV 863006.612p 0.563673mV 863009.57p 0.563673mV 864018.723p 0.603491mV 864036.727p 0.638979mV 865001.803p 0.551358mV 865020.915p 0.586293mV 865021.692p 0.586293mV 865033.655p 0.551099mV 865070.167p 0.585999mV 865076.925p 0.603544mV 865082.502p 0.585979mV 865083.989p 0.585979mV 865114.421p 0.62127mV 865132.271p 0.586533mV 865141.485p 0.586832mV 865146.607p 0.569457mV 865147.461p 0.569457mV 865157.652p 0.604893mV 866003.597p 0.553537mV 866020.208p 0.553336mV 866070.786p 0.658946mV 867007.593p 0.565666mV 867018.148p 0.530531mV 867043.618p 0.51284mV 867048.349p 0.530322mV 867075.992p 0.564863mV 867140.804p 0.581223mV 867145.195p 0.563574mV 867190.645p 0.545229mV 867207.89p 0.527381mV 867210.556p 0.509701mV 867220.077p 0.474323mV 868026.689p 0.532812mV 868032.921p 0.515277mV 868078.109p 0.462086mV 869004.985p 0.550432mV 869018.159p 0.532792mV 869032.612p 0.550231mV 869055.594p 0.532319mV 869076.547p 0.602014mV 869082.564p 0.619444mV 869101.546p 0.619165mV 869113.866p 0.619162mV 869114.627p 0.619162mV 869122.765p 0.619249mV 869132.144p 0.654507mV 869135.736p 0.672157mV 870009.19p 0.563807mV 870021.947p 0.58121mV 870031.369p 0.581157mV 870051.954p 0.546093mV 870061.761p 0.546144mV 870068.196p 0.563736mV 870112.435p 0.511163mV 870121.54p 0.546195mV 870131.009p 0.546077mV 871028.54p 0.533419mV 871088.532p 0.498374mV 871088.861p 0.498374mV 871094.043p 0.480726mV 871097.435p 0.463067mV 872006.55p 0.530564mV 872014.339p 0.513045mV 872053.071p 0.547878mV 872076.096p 0.564867mV 872095.585p 0.56441mV 872101.246p 0.581836mV 872141.471p 0.580759mV 872141.591p 0.580759mV 872171.814p 0.685157mV 872200.59p 0.650032mV 872205.886p 0.667668mV 872208.881p 0.667668mV 872231.91p 0.615802mV 872236.9p 0.598503mV 873029.145p 0.531811mV 873050.135p 0.51437mV 873055.438p 0.531946mV 873056.259p 0.531946mV 873063.661p 0.514387mV 873081.164p 0.514282mV 873087.264p 0.531769mV 873089.695p 0.531769mV 873140.915p 0.512615mV 873144.188p 0.512615mV 874002.234p 0.547469mV 874015.503p 0.565114mV 874042.141p 0.547968mV 874042.803p 0.547968mV 874086.738p 0.566563mV 874104.348p 0.549427mV 874104.355p 0.549427mV 874118.295p 0.567522mV 874124.749p 0.585249mV 875013.595p 0.518834mV 875036.994p 0.501053mV 876023.36p 0.581218mV 877037.622p 0.570876mV 877045.342p 0.605919mV 877049.16p 0.605919mV 877052.5p 0.623457mV 877053.666p 0.623457mV 877115.243p 0.571706mV 877127.805p 0.572002mV 877163.805p 0.555958mV 878018.815p 0.536172mV 878024.77p 0.553747mV 878027.724p 0.571317mV 878075.03p 0.571652mV 878154.719p 0.589983mV 878166.467p 0.572558mV 878177.822p 0.537611mV 878187.736p 0.572922mV 878214.036p 0.556195mV 879046.364p 0.463293mV 879055.05p 0.498331mV 880004.749p 0.550896mV 880011.863p 0.515739mV 880022.057p 0.515671mV 880023.032p 0.515671mV 880029.554p 0.498062mV 880062.15p 0.514614mV 881004.316p 0.549043mV 881050.81p 0.514455mV 882043.287p 0.511981mV 882053.855p 0.51205mV 882074.689p 0.476982mV 882087.507p 0.49443mV 883017.894p 0.569783mV 883041.912p 0.551992mV 883128.994p 0.533083mV 884008.233p 0.570931mV 884014.509p 0.553381mV 884032.397p 0.553451mV 884054.143p 0.553513mV 884081.736p 0.588866mV 884130.503p 0.625088mV 885037.959p 0.500064mV 885072.282p 0.552066mV 885077.015p 0.53439mV 886006.93p 0.530247mV 886031.444p 0.512812mV 886038.777p 0.530376mV 886039.431p 0.530376mV 886051.513p 0.512759mV 886064.695p 0.547759mV 886070.408p 0.582728mV 886085.19p 0.565026mV 886100.257p 0.617688mV 886103.46p 0.617688mV 887013.038p 0.552737mV 887021.518p 0.517666mV 887049.558p 0.499989mV 888005.815p 0.530047mV 889017.784p 0.528861mV 889040.525p 0.511061mV 889045.374p 0.528518mV 889068.572p 0.563126mV 889104.719p 0.579833mV 889135.084p 0.526443mV 889159.707p 0.560951mV 889180.173p 0.612432mV 889183.351p 0.612432mV 889202.071p 0.611508mV 889218.465p 0.628408mV 890003.531p 0.554222mV 890028.133p 0.536402mV 890051.618p 0.55348mV 890070.342p 0.552998mV 890072.788p 0.552998mV 890084.773p 0.552697mV 890088.21p 0.535mV 890101.876p 0.587068mV 890127.593p 0.638735mV 890142.709p 0.65594mV 890166.016p 0.708483mV 890174.394p 0.69098mV 890178.516p 0.673525mV 891016.143p 0.570165mV 891019.608p 0.570165mV 891046.801p 0.569905mV 891049.417p 0.569905mV 891074.992p 0.552179mV 891106.642p 0.604779mV 891110.186p 0.58725mV 891111.291p 0.58725mV 891129.363p 0.604994mV 891142.49p 0.62286mV 891171.358p 0.519011mV 891184.825p 0.519495mV 891212.539p 0.520931mV 892039.084p 0.570043mV 892053.714p 0.5525mV 892067.876p 0.535023mV 892071.146p 0.51749mV 892074.42p 0.51749mV 892106.062p 0.429459mV 893004.507p 0.547005mV 893017.695p 0.564502mV 893033.335p 0.546928mV 893065.256p 0.529318mV 893083.683p 0.511558mV 893108.98p 0.563736mV 893113.068p 0.546078mV 893115.126p 0.528422mV 893115.555p 0.528422mV 894001.076p 0.552885mV 894009.642p 0.570461mV 894026.4p 0.570589mV 895013.479p 0.582443mV 895018.339p 0.600015mV 895022.957p 0.617601mV 895029.135p 0.635204mV 895039.878p 0.635372mV 896003.95p 0.548044mV 896022.533p 0.548038mV 896048.87p 0.635989mV 896064.489p 0.618779mV 896069.478p 0.601439mV 897021.34p 0.581466mV 897025.066p 0.564mV 897025.479p 0.564mV 897033.296p 0.581659mV 897055.861p 0.599959mV 897059.93p 0.599959mV 898024.871p 0.550974mV 898044.712p 0.550954mV 899012.67p 0.518717mV 899020.866p 0.553797mV 899044.788p 0.588796mV 899057.976p 0.606352mV 899058.812p 0.606352mV 899060.659p 0.623944mV 899074.867p 0.62407mV 899081.137p 0.624318mV 899090.728p 0.624658mV 899091.19p 0.624658mV 900014.053p 0.584727mV 901007.04p 0.569478mV 901011.732p 0.587027mV 901037.113p 0.639848mV 902002.393p 0.548757mV 902005.483p 0.566264mV 902012.808p 0.548655mV 902012.919p 0.548655mV 902031.421p 0.583635mV 902032.621p 0.583635mV 902069.639p 0.601599mV 902074.353p 0.619307mV 902076.816p 0.601966mV 903007.656p 0.53431mV 903017.929p 0.499243mV 903018.05p 0.499243mV 903023.369p 0.516813mV 903038.44p 0.499171mV 903045.222p 0.499005mV 903066.044p 0.568634mV 903093.855p 0.515226mV 903103.067p 0.514882mV 904015.529p 0.563409mV 904047.839p 0.493208mV 904073.075p 0.510487mV 904096.764p 0.527209mV 904101.125p 0.54449mV 905006.007p 0.564mV 905017.884p 0.528958mV 905024.897p 0.51144mV 905056.529p 0.494mV 905099.365p 0.528737mV 905122.539p 0.545863mV 905130.36p 0.545659mV 906013.69p 0.551366mV 906015.55p 0.568896mV 906019.564p 0.568896mV 906038.256p 0.568819mV 906046.458p 0.603928mV 906056.901p 0.603966mV 906079.139p 0.569112mV 906082.406p 0.551655mV 906095.117p 0.569517mV 906110.064p 0.517185mV 906137.514p 0.535261mV 906138.687p 0.535261mV 906139.029p 0.535261mV 906165.011p 0.606293mV 906165.508p 0.606293mV 907010.773p 0.511791mV 907028.844p 0.564379mV 907034.899p 0.546777mV 907044.106p 0.5467mV 907139.722p 0.597442mV 907148.446p 0.632448mV 907158.26p 0.667519mV 908023.487p 0.58672mV 908043.291p 0.551744mV 908044.668p 0.551744mV 908066.625p 0.534298mV 908129.868p 0.533298mV 908148.691p 0.497537mV 909003.998p 0.546335mV 909016.791p 0.528827mV 909051.197p 0.546381mV 909072.985p 0.581424mV 909079.051p 0.598966mV 909107.638p 0.599339mV 910013.845p 0.51759mV 910018.041p 0.535109mV 910031.399p 0.552475mV 910083.835p 0.516202mV 910088.276p 0.498465mV 911029.489p 0.605348mV 911037.244p 0.60538mV 911078.014p 0.53607mV 911078.078p 0.53607mV 911092.241p 0.483975mV 911163.952p 0.484398mV 911175.996p 0.466635mV 911188.575p 0.501493mV 911236.174p 0.569778mV 911286.397p 0.637701mV 911303.332p 0.584576mV 911306.651p 0.601959mV 911339.393p 0.636105mV 911348.215p 0.600728mV 911351.001p 0.618137mV 911354.623p 0.618137mV 911372.132p 0.652626mV 911402.729p 0.651875mV 911424.665p 0.616468mV 911456.563p 0.66834mV 911466.346p 0.703216mV 911489.249p 0.702972mV 911506.094p 0.632798mV 912016.443p 0.529426mV 912017.805p 0.529426mV 912074.965p 0.582364mV 912084.955p 0.582635mV 912095.657p 0.53055mV 912100.194p 0.548278mV 912119.913p 0.531366mV 912126.191p 0.566835mV 912129.117p 0.566835mV 913008.595p 0.563827mV 913049.225p 0.492982mV 914013.838p 0.517417mV 914014.842p 0.517417mV 914026.526p 0.499647mV 914043.032p 0.551895mV 914066.799p 0.60369mV 914074.737p 0.621108mV 914089.453p 0.638375mV 914089.914p 0.638375mV 914094.274p 0.655877mV 914112.413p 0.655927mV 915006.855p 0.534089mV 915013.503p 0.51654mV 915035.964p 0.463743mV 915046.02p 0.463557mV 915049.869p 0.463557mV 916019.059p 0.570139mV 916045.461p 0.605413mV 916057.73p 0.605578mV 917003.728p 0.553881mV 917037.258p 0.571304mV 917047.02p 0.60636mV 917061.821p 0.623937mV 917077.715p 0.571476mV 917093.368p 0.58939mV 917094.953p 0.58939mV 917117.446p 0.537706mV 918012.858p 0.511336mV 918012.966p 0.511336mV 918016.246p 0.49378mV 918054.594p 0.475796mV 919000.463p 0.548514mV 919011.123p 0.583733mV 919012.621p 0.583733mV 919022.94p 0.583864mV 920000.487p 0.554335mV 920016.203p 0.60713mV 920033.57p 0.624921mV 920035.428p 0.607498mV 921028.22p 0.637108mV 921039.681p 0.63718mV 922009.693p 0.535934mV 922034.8p 0.482861mV 923044.845p 0.652991mV 923047.596p 0.635512mV 923051.522p 0.653176mV 923059.135p 0.635775mV 924008.153p 0.569322mV 924010.381p 0.586897mV 924036.427p 0.67497mV 924040.502p 0.657554mV 925014.194p 0.550685mV 925037.283p 0.568271mV 925076.899p 0.53347mV 925085.97p 0.568624mV 925088.846p 0.568624mV 925095.594p 0.568666mV 925105.617p 0.568734mV 925124.202p 0.586456mV 925132.019p 0.621763mV 926024.539p 0.588913mV 926026.28p 0.571428mV 926027.032p 0.571428mV 926077.185p 0.53755mV 926091.904p 0.520345mV 926094.051p 0.520345mV 926161.456p 0.557346mV 927031.352p 0.621404mV 927044.464p 0.621456mV 927049.033p 0.603973mV 928018.231p 0.598346mV 928018.244p 0.598346mV 928020.523p 0.615927mV 929001.251p 0.546548mV 929008.866p 0.564086mV 930016.281p 0.499378mV 930019.706p 0.499378mV 930020.73p 0.481803mV 930023.819p 0.481803mV 930036.978p 0.499167mV 930086.041p 0.532383mV 931020.885p 0.548143mV 931025.697p 0.530591mV 931034.679p 0.54816mV 931044.546p 0.583284mV 931046.676p 0.600853mV 931054.966p 0.583315mV 931063.07p 0.583419mV 931075.691p 0.53105mV 931080.111p 0.548712mV 931088.993p 0.566371mV 931105.602p 0.566902mV 931116.227p 0.532227mV 931116.648p 0.532227mV 931117.325p 0.532227mV 932013.026p 0.586619mV 933026.181p 0.642301mV 933030.919p 0.624868mV 934002.073p 0.551228mV 934013.863p 0.586444mV 934015.408p 0.568941mV 934033.501p 0.551615mV 934045.343p 0.604556mV 934047.381p 0.604556mV 935004.44p 0.554007mV 935012.812p 0.553962mV 935028.214p 0.606564mV 935089.541p 0.572236mV 935092.066p 0.5899mV 935109.394p 0.642935mV 935110.218p 0.625574mV 936001.793p 0.545928mV 936034.075p 0.54583mV 936067.213p 0.528034mV 936086.527p 0.562806mV 936100.138p 0.544945mV 936137.062p 0.631693mV 936162.115p 0.578605mV 936165.287p 0.560992mV 936181.297p 0.613481mV 936188.128p 0.595862mV 936231.252p 0.612892mV 936262.844p 0.542192mV 936264.428p 0.542192mV 936265.592p 0.559644mV 936272.421p 0.577065mV 936299.013p 0.628911mV 936321.376p 0.610638mV 936330.129p 0.575278mV 936337.799p 0.592677mV 936362.07p 0.644273mV 936392.588p 0.642962mV 936394.261p 0.642962mV 936400.74p 0.677637mV 936418.551p 0.659513mV 936451.333p 0.710682mV 936470.699p 0.67487mV 937011.698p 0.546748mV 937018.288p 0.564303mV 937019.407p 0.564303mV 937030.464p 0.581876mV 937043.967p 0.581937mV 937070.932p 0.547246mV 937086.018p 0.60023mV 937099.534p 0.600512mV 937106.289p 0.600873mV 937108.239p 0.600873mV 938035.223p 0.599621mV 938055.808p 0.565075mV 938058.501p 0.565075mV 938095.874p 0.496692mV 938121.433p 0.480395mV 938126.733p 0.463123mV 938133.956p 0.480873mV 939002.44p 0.550579mV 939004.536p 0.550579mV 939052.46p 0.65579mV 939060.893p 0.656005mV 939065.103p 0.673687mV 940016.098p 0.500687mV 940038.902p 0.500233mV 941009.1p 0.570252mV 941024.786p 0.587674mV 942023.369p 0.51339mV 942044.723p 0.443153mV 943069.199p 0.642533mV 944010.518p 0.586812mV 944012.439p 0.586812mV 944023.459p 0.622024mV 944026.088p 0.639652mV 944036.764p 0.604782mV 944051.586p 0.587835mV 946031.688p 0.512881mV 946032.577p 0.512881mV 946033.245p 0.512881mV 946048.399p 0.460103mV 946057.768p 0.495024mV 946073.02p 0.51205mV 947016.759p 0.49431mV 947039.063p 0.528962mV 947042.789p 0.54635mV 947047.018p 0.563722mV 947048.391p 0.563722mV 947070.04p 0.580456mV 947088.096p 0.597618mV 947098.502p 0.56231mV 948010.533p 0.512752mV 948022.083p 0.512668mV 948056.261p 0.494197mV 948060.019p 0.511506mV 949042.935p 0.5514mV 949054.825p 0.516071mV 949058.431p 0.498399mV 950034.762p 0.588094mV 951026.752p 0.566253mV 951031.877p 0.54864mV 951043.491p 0.583659mV 951093.745p 0.61911mV 952013.394p 0.55072mV 952019.622p 0.533149mV 952103.889p 0.583536mV 952121.691p 0.617912mV 952121.752p 0.617912mV 952121.943p 0.617912mV 952148.76p 0.634847mV 952149.481p 0.634847mV 952158.163p 0.59959mV 952160.811p 0.581974mV 952181.061p 0.616828mV 952203.87p 0.686854mV 952217.483p 0.669361mV 952229.439p 0.669515mV 952281.971p 0.548833mV 952294.006p 0.584278mV 952301.287p 0.584648mV 952324.002p 0.585511mV 953028.445p 0.598988mV 953036.603p 0.634167mV 953058.871p 0.599509mV 954008.359p 0.536211mV 954015.403p 0.53611mV 954038.503p 0.606023mV 954064.01p 0.62346mV 954072.405p 0.623531mV 954078.781p 0.606054mV 954086.234p 0.571189mV 954096.064p 0.571476mV 955000.921p 0.546894mV 955002.567p 0.546894mV 955018.504p 0.564495mV 955047.499p 0.599816mV 955064.39p 0.617644mV 956005.283p 0.536573mV 956089.834p 0.571253mV 956093.291p 0.588771mV 956095.298p 0.571175mV 956106.654p 0.571131mV 956124.842p 0.588642mV 956148.017p 0.641544mV 957001.863p 0.548348mV 957046.1p 0.460012mV 958021.182p 0.546889mV 958022.686p 0.546889mV 958039.391p 0.529398mV 958039.79p 0.529398mV 958046.598p 0.529431mV 958109.439p 0.528454mV 958121.486p 0.51032mV 959002.877p 0.553993mV 959048.749p 0.53666mV 959049.77p 0.53666mV 959053.183p 0.554208mV 959057.753p 0.536629mV 959058.343p 0.536629mV 959058.937p 0.536629mV 959082.028p 0.518938mV 959090.815p 0.553911mV 959104.137p 0.51863mV 959105.702p 0.536093mV 959125.938p 0.535586mV 959144.721p 0.517565mV 959146.042p 0.499839mV 960014.199p 0.549876mV 960014.393p 0.549876mV 960033.416p 0.549679mV 960036.89p 0.567164mV 960071.509p 0.584485mV 960074.554p 0.584485mV 960082.128p 0.549438mV 960104.543p 0.549599mV 960108.337p 0.567198mV 960135.41p 0.497149mV 960170.419p 0.549361mV 960171.543p 0.549361mV 960185.68p 0.566616mV 960197.151p 0.566415mV 960197.695p 0.566415mV 960209.984p 0.566236mV 961005.669p 0.570907mV 961027.346p 0.536039mV 961066.414p 0.465891mV 961081.74p 0.447927mV 962069.276p 0.529688mV 962075.753p 0.564439mV 962081.34p 0.546727mV 962115.749p 0.598091mV 962118.169p 0.598091mV 962130.733p 0.615137mV 962141.684p 0.64992mV 962150.17p 0.649695mV 962169.535p 0.702227mV 962170.186p 0.719798mV 963040.783p 0.586861mV 963045.538p 0.604462mV 964009.483p 0.534788mV 964018.566p 0.534711mV 964051.364p 0.516558mV 964083.753p 0.55048mV 964086.913p 0.567764mV 965015.42p 0.534831mV 965019.753p 0.534831mV 965021.951p 0.517318mV 966028.948p 0.606492mV 966030.124p 0.588941mV 966044.26p 0.589021mV 966081.012p 0.624929mV 967030.139p 0.546107mV 967076.82p 0.563672mV 967115.859p 0.599333mV 968040.116p 0.588328mV 969000.304p 0.553374mV 969028.268p 0.500789mV 970005.043p 0.563044mV 970016.147p 0.598059mV 970049.903p 0.562912mV 970101.68p 0.51002mV 970102.826p 0.51002mV 970114.199p 0.509788mV 971010.978p 0.547889mV 971023.953p 0.512842mV 971057.67p 0.49532mV 971123.467p 0.510958mV 972033.607p 0.655809mV 972037.096p 0.673445mV 972037.784p 0.673445mV 973057.32p 0.458878mV 974032.314p 0.58461mV 974040.632p 0.584726mV 975021.682p 0.588071mV 975048.191p 0.500545mV 975102.434p 0.482516mV 976033.636p 0.512089mV 976062.295p 0.441426mV 977002.478p 0.551193mV 977023.975p 0.586349mV 977048.813p 0.639252mV 977064.217p 0.692231mV 977064.358p 0.692231mV 978027.149p 0.601894mV 978031.937p 0.619474mV 979012.68p 0.512492mV 979023.802p 0.547677mV 979032.24p 0.512595mV 979035.284p 0.530169mV 979045.424p 0.49504mV 979053.571p 0.477459mV 979056.004p 0.49498mV 979092.522p 0.511702mV 980006.502p 0.535381mV 980009.849p 0.535381mV 980019.432p 0.500206mV 980025.127p 0.500099mV 980040.743p 0.48221mV 980044.022p 0.48221mV 980044.743p 0.48221mV 981001.328p 0.549203mV 981015.609p 0.531826mV 981015.974p 0.531826mV 981020.225p 0.54945mV 981046.571p 0.602511mV 982013.538p 0.548914mV 982017.601p 0.566467mV 982019.935p 0.566467mV 982022.3p 0.58402mV 982056.601p 0.637143mV 982062.108p 0.654842mV 983051.062p 0.621451mV 983078.455p 0.674134mV 983083.908p 0.69176mV 984032.981p 0.586319mV 984035.402p 0.568826mV 984053.902p 0.551541mV 984086.977p 0.56993mV 984090.109p 0.587604mV 984095.342p 0.570196mV 985027.004p 0.535263mV 985035.39p 0.535302mV 985064.962p 0.482629mV 985073.788p 0.447419mV 986039.521p 0.497192mV 986046.532p 0.497125mV 986064.434p 0.514404mV 986069.027p 0.496725mV 986070.755p 0.479039mV 987006.524p 0.528864mV 987011.448p 0.546405mV 987024.103p 0.546352mV 987042.26p 0.546267mV 987046.313p 0.528675mV 987075.825p 0.598657mV 987097.519p 0.598684mV 987113.41p 0.581418mV 987126.925p 0.599403mV 988000.048p 0.546335mV 988013.6p 0.581488mV 989000.456p 0.553398mV 989030.559p 0.517868mV 989041.218p 0.482536mV 989057.827p 0.499574mV 990014.337p 0.514992mV 990021.331p 0.514985mV 990064.403p 0.549431mV 990085.204p 0.601259mV 990105.04p 0.565582mV 990108.321p 0.565582mV 991007.171p 0.535453mV 991021.266p 0.482701mV 991021.677p 0.482701mV 992009.545p 0.532702mV 992028.723p 0.497472mV 992030.618p 0.479859mV 992047.211p 0.532205mV 992051.469p 0.549598mV 992062.071p 0.549274mV 993000.973p 0.548525mV 993012.94p 0.583726mV 993026.516p 0.56635mV 993049.245p 0.566773mV 993056.187p 0.60215mV 994009.647p 0.564639mV 994039.866p 0.600074mV 995033.742p 0.622261mV 996015.425p 0.532573mV 996053.6p 0.584524mV 996061.247p 0.5843mV 997002.05p 0.548792mV 997006.399p 0.531201mV 997009.691p 0.531201mV 997043.567p 0.583644mV 998004.193p 0.550237mV 998035.089p 0.497727mV 998046.851p 0.462594mV 998051.185p 0.444995mV 998058.094p 0.462487mV 998072.522p 0.479616mV 998073.931p 0.479616mV 999000.628p 0.546427mV 999021.397p 0.546648mV 999034.182p 0.581894mV 999058.936p 0.564868mV 999063.619p 0.582553mV 999071.763p 0.582871mV 999076.932p 0.565523mV)
.ENDS conductors__anyBias-Lk_0_702

.SUBCKT conductors__anyBias-Lk_0_703 bottom out
VrampSppl@0 bottom out pwl (0 0 2.626p 0.587029mV 9.16p 0.586807mV 1010.55p 0.55707mV 2003.011p 0.521306mV 2017.865p 0.516222mV 2049.239p 0.55777mV 2063.421p 0.593515mV 2134.38p 0.396969mV 3004.63p 0.497197mV 3009.668p 0.497386mV 3015.246p 0.503059mV 3021.227p 0.508584mV 3036.491p 0.548743mV 3056.112p 0.618275mV 3078.865p 0.743433mV 4006.61p 0.598003mV 4014.536p 0.591409mV 4018.973p 0.591413mV 4024.43p 0.597974mV 4044.994p 0.665216mV 4050.965p 0.727128mV 4059.298p 0.756222mV 5001.999p 0.531085mV 5002.467p 0.531085mV 5038.347p 0.502136mV 5094.791p 0.616952mV 5122.937p 0.775054mV 6044.332p 0.549192mV 6047.645p 0.56125mV 6047.803p 0.56125mV 6050.245p 0.579605mV 6076.369p 0.719057mV 6078.354p 0.719057mV 6078.879p 0.719057mV 7025.438p 0.644216mV 7040.383p 0.677427mV 7044.48p 0.677427mV 7053.015p 0.680161mV 7055.518p 0.685877mV 7058.78p 0.685877mV 7065.342p 0.693548mV 7078.81p 0.692203mV 7081.941p 0.683541mV 7086.85p 0.669533mV 7087.971p 0.669533mV 7091.535p 0.662609mV 8001.572p 0.517914mV 8062.014p 0.472462mV 8079.816p 0.492149mV 8088.444p 0.526239mV 8097.905p 0.571848mV 8103.15p 0.597745mV 8134.259p 0.76826mV 8134.334p 0.76826mV 9017.605p 0.533638mV 9028.063p 0.502626mV 9041.972p 0.46382mV 10015.957p 0.527407mV 11025.849p 0.561189mV 11049.928p 0.500682mV 12015.671p 0.587781mV 13019.122p 0.560125mV 13050.9p 0.602324mV 13075.503p 0.701708mV 13090.788p 0.717783mV 13103.647p 0.739845mV 14004.679p 0.597016mV 14021.903p 0.586259mV 14034.508p 0.595061mV 14053.919p 0.628443mV 14064.579p 0.666317mV 14073.376p 0.694068mV 14085.638p 0.732771mV 14090.627p 0.747729mV 14091.777p 0.747729mV 14095.232p 0.757631mV 14097.682p 0.757631mV 15013.802p 0.566755mV 15019.42p 0.566503mV 15027.574p 0.585217mV 15056.121p 0.647816mV 15056.909p 0.647816mV 15074.853p 0.695582mV 15083.609p 0.737442mV 15086.074p 0.769182mV 15086.456p 0.769182mV 15089.995p 0.769182mV 16004.96p 0.51732mV 16056.86p 0.605226mV 16059.189p 0.605226mV 16074.697p 0.673323mV 16082.326p 0.71547mV 17042.248p 0.456206mV 17071.667p 0.35704mV 18028.91p 0.600848mV 18049.831p 0.669079mV 18060.546p 0.679625mV 18061.709p 0.679625mV 18079.839p 0.703727mV 18096.027p 0.753146mV 19008.371p 0.51628mV 19038.32p 0.567799mV 19085.732p 0.71399mV 19089.309p 0.71399mV 20008.652p 0.570178mV 20011.427p 0.576764mV 20013.896p 0.576764mV 20019.006p 0.589779mV 20027.76p 0.622698mV 20048.291p 0.680891mV 20057.526p 0.732662mV 21042.875p 0.554465mV 21043.024p 0.554465mV 21049.596p 0.553923mV 21051.64p 0.547108mV 21075.49p 0.44264mV 22001.265p 0.540201mV 22032.142p 0.569784mV 22058.057p 0.608576mV 22082.459p 0.700263mV 22101.712p 0.685649mV 22116.298p 0.618753mV 22116.901p 0.618753mV 22131.655p 0.538357mV 22138.949p 0.499441mV 23024.938p 0.518236mV 23059.659p 0.551722mV 23063.413p 0.568402mV 23068.699p 0.591394mV 23080.343p 0.6364mV 23101.495p 0.774477mV 24000.06p 0.51361mV 24014.375p 0.505297mV 24016.603p 0.491345mV 24033.823p 0.40966mV 25029.011p 0.528913mV 25029.262p 0.528913mV 25051.705p 0.520604mV 25121.929p 0.564949mV 25143.025p 0.68669mV 25144.416p 0.68669mV 25149.378p 0.721319mV 26021.134p 0.522922mV 26041.447p 0.492833mV 26056.037p 0.479646mV 26057.824p 0.479646mV 26084.597p 0.491478mV 27021.006p 0.547717mV 27042.395p 0.50122mV 27045.266p 0.476666mV 27046.107p 0.476666mV 28012.779p 0.583398mV 28048.699p 0.557003mV 28052.812p 0.539347mV 28054.928p 0.539347mV 29002.118p 0.574701mV 29007.265p 0.573688mV 30002.869p 0.584658mV 30035.466p 0.53546mV 30035.892p 0.53546mV 30043.161p 0.517916mV 30060.19p 0.471024mV 30120.104p 0.540192mV 30120.259p 0.540192mV 30132.874p 0.59478mV 30143.59p 0.63724mV 30160.231p 0.7535mV 31001.235p 0.573898mV 31041.854p 0.555904mV 31119.772p 0.380679mV 32012.035p 0.504304mV 32014.166p 0.504304mV 32026.036p 0.517795mV 32040.276p 0.52271mV 32095.051p 0.697382mV 32101.044p 0.72804mV 32108.998p 0.76585mV 33026.303p 0.537021mV 33039.775p 0.533435mV 33048.205p 0.529437mV 33065.111p 0.507128mV 33094.759p 0.600258mV 33114.522p 0.727113mV 33114.993p 0.727113mV 33118.721p 0.766787mV 34004.228p 0.498021mV 34025.182p 0.49434mV 34033.541p 0.498837mV 34040.723p 0.513097mV 34069.922p 0.522317mV 34070.308p 0.52485mV 34114.893p 0.409817mV 34130.194p 0.361814mV 34150.38p 0.345335mV 34204.542p 0.496731mV 34227.831p 0.590591mV 34240.074p 0.624643mV 34257.635p 0.656167mV 35013.496p 0.55139mV 35019.106p 0.538114mV 35037.008p 0.496985mV 35089.968p 0.345132mV 36022.898p 0.547711mV 36040.848p 0.616716mV 36053.251p 0.633675mV 36060.662p 0.652563mV 36069.543p 0.666008mV 37007.03p 0.507812mV 37009.256p 0.507812mV 37044.084p 0.571596mV 37047.901p 0.583987mV 37048.302p 0.583987mV 37060.734p 0.647529mV 37069.015p 0.673679mV 37073.963p 0.694167mV 37080.915p 0.756337mV 38012.176p 0.507072mV 38062.819p 0.615292mV 38085.608p 0.714448mV 38091.116p 0.737627mV 38097.518p 0.76805mV 39015.423p 0.57945mV 39021.575p 0.586328mV 39035.858p 0.583014mV 39068.419p 0.551032mV 39069.148p 0.551032mV 39103.989p 0.492326mV 39124.361p 0.420402mV 39165.943p 0.35509mV 40002.868p 0.58433mV 40005.3p 0.583525mV 40011.987p 0.589234mV 40036.811p 0.551826mV 40044.462p 0.546065mV 40051.635p 0.553446mV 40061.457p 0.560781mV 40070.311p 0.555653mV 40096.77p 0.508902mV 40120.451p 0.451609mV 40192.462p 0.563073mV 40195.02p 0.568247mV 40213.623p 0.584356mV 40219.332p 0.589978mV 40244.489p 0.603403mV 40248.5p 0.610891mV 40275.243p 0.709621mV 40285.408p 0.765137mV 41040.551p 0.577557mV 41097.412p 0.682874mV 42017.572p 0.625574mV 42046.656p 0.741133mV 43012.086p 0.50806mV 43022.723p 0.501203mV 43030.309p 0.505833mV 43065.114p 0.445386mV 43126.216p 0.397833mV 43130.929p 0.400737mV 43160.998p 0.442776mV 43168.901p 0.458424mV 43194.968p 0.585453mV 44030.358p 0.632159mV 44067.084p 0.760033mV 45006.97p 0.508078mV 45055.229p 0.374576mV 46032.657p 0.569709mV 46034.932p 0.569709mV 46049.725p 0.588824mV 46067.596p 0.642587mV 46087.232p 0.704633mV 47072.714p 0.525531mV 48031.919p 0.414496mV 48035.969p 0.398562mV 49016.845p 0.50959mV 49040.712p 0.460935mV 49055.766p 0.446415mV 50004.009p 0.519927mV 50004.933p 0.519927mV 50012.63p 0.52613mV 50025.633p 0.543652mV 50060.725p 0.486974mV 50092.463p 0.476578mV 50101.646p 0.498941mV 50105.433p 0.518913mV 50112.086p 0.53227mV 50117.571p 0.55173mV 50173.908p 0.767016mV 50179.114p 0.769817mV 50181.3p 0.767817mV 50184.17p 0.767817mV 50191.333p 0.761776mV 50192.87p 0.761776mV 50203.059p 0.773378mV 51008.018p 0.497058mV 51008.699p 0.497058mV 51008.959p 0.497058mV 51024.496p 0.492779mV 51056.986p 0.514033mV 51094.492p 0.579724mV 51107.133p 0.609728mV 51129.393p 0.645864mV 51171.75p 0.705345mV 51175.182p 0.72189mV 51175.981p 0.72189mV 52008.66p 0.555281mV 52050.544p 0.495918mV 52053.788p 0.495918mV 52055.361p 0.482203mV 53005.54p 0.600163mV 53012.121p 0.606313mV 53012.901p 0.606313mV 53030.575p 0.634599mV 54013.121p 0.5335mV 54014.461p 0.5335mV 54020.476p 0.541285mV 54024.347p 0.541285mV 54039.491p 0.587083mV 54044.361p 0.6067mV 54050.905p 0.62787mV 54073.216p 0.72625mV 55000.05p 0.531964mV 56048.527p 0.506755mV 56075.42p 0.458897mV 56106.871p 0.417785mV 56126.505p 0.363627mV 56126.737p 0.363627mV 57023.364p 0.605004mV 57034.718p 0.652036mV 57064.634p 0.707814mV 57075.038p 0.763148mV 58017.161p 0.570465mV 58041.767p 0.520003mV 58050.077p 0.503396mV 58069.352p 0.511176mV 58125.375p 0.383561mV 59024.404p 0.544053mV 59055.604p 0.447723mV 59065.605p 0.412513mV 59085.704p 0.332422mV 60076.008p 0.532184mV 60082.382p 0.538681mV 60096.738p 0.595508mV 60108.896p 0.652804mV 61008.257p 0.583851mV 61024.616p 0.585461mV 61044.189p 0.615925mV 61061.717p 0.640028mV 61073.323p 0.63026mV 61117.355p 0.527828mV 61168.331p 0.485141mV 62041.733p 0.569964mV 62053.415p 0.587287mV 62083.997p 0.671401mV 62092.182p 0.683161mV 62101.083p 0.685578mV 62108.829p 0.691187mV 62120.89p 0.713333mV 62129.086p 0.710213mV 63049.498p 0.523312mV 63051.604p 0.528546mV 63065.959p 0.53073mV 63125.444p 0.464574mV 63135.93p 0.424996mV 63151.901p 0.35719mV 64023.271p 0.538288mV 64054.166p 0.402552mV 65022.833p 0.518425mV 65023.382p 0.518425mV 66001.88p 0.575779mV 66006.365p 0.575982mV 66029.313p 0.515241mV 66061.282p 0.410724mV 66074.41p 0.409857mV 66092.006p 0.397632mV 66103.921p 0.348855mV 67015.696p 0.492345mV 67024.871p 0.473373mV 67032.489p 0.453088mV 67046.204p 0.390117mV 68034.399p 0.47084mV 68036.284p 0.445705mV 69007.335p 0.603521mV 69024.993p 0.607387mV 69030.709p 0.60555mV 69067.389p 0.601088mV 69079.696p 0.568012mV 69084.978p 0.542427mV 69092.006p 0.497733mV 69094.533p 0.497733mV 69127.989p 0.367923mV 70004.982p 0.580999mV 70006.113p 0.580315mV 70008.665p 0.580315mV 70011.685p 0.586126mV 70012.842p 0.586126mV 70033.934p 0.611779mV 70054.299p 0.668464mV 70057.736p 0.683978mV 71002.332p 0.553204mV 71026.348p 0.544885mV 72010.185p 0.523571mV 72016.131p 0.522174mV 72046.763p 0.542035mV 72058.429p 0.543744mV 72070.057p 0.574423mV 72075.882p 0.597279mV 72088.855p 0.649899mV 73035.599p 0.518172mV 73037.405p 0.518172mV 73085.525p 0.439733mV 73117.214p 0.453293mV 73154.62p 0.564888mV 73163.481p 0.560294mV 73193.819p 0.58658mV 73205.746p 0.624053mV 74009.88p 0.522004mV 75012.498p 0.523073mV 75061.563p 0.50552mV 75101.288p 0.464458mV 75147.848p 0.461286mV 75198.437p 0.694338mV 75207.407p 0.731931mV 76025.845p 0.618361mV 76044.849p 0.583894mV 76076.881p 0.47634mV 76109.624p 0.515883mV 76170.198p 0.562919mV 76182.473p 0.55266mV 76195.166p 0.553393mV 76204.421p 0.545277mV 76230.67p 0.603756mV 76253.536p 0.688545mV 76258.175p 0.726782mV 76260.016p 0.759635mV 77027.655p 0.585227mV 77062.292p 0.471765mV 77076.039p 0.417746mV 78059.644p 0.757333mV 79029.742p 0.605746mV 79048.095p 0.615144mV 79049.693p 0.615144mV 79053.975p 0.624679mV 79091.491p 0.770088mV 79092.045p 0.770088mV 80003.236p 0.497538mV 80060.113p 0.661749mV 81030.733p 0.504016mV 81031.582p 0.504016mV 81040.937p 0.507962mV 81070.739p 0.512735mV 81075.419p 0.509336mV 81136.403p 0.50174mV 81161.696p 0.512444mV 81167.002p 0.51758mV 81168.367p 0.51758mV 81170.223p 0.516181mV 81187.219p 0.548553mV 81208.417p 0.590641mV 81222.752p 0.642755mV 81226.123p 0.648418mV 81229.015p 0.648418mV 81235.541p 0.655255mV 81237.224p 0.655255mV 81247.213p 0.664608mV 81251.234p 0.667153mV 81287.754p 0.758386mV 82024.89p 0.576041mV 82050.039p 0.615971mV 82070.269p 0.616007mV 82075.524p 0.620217mV 82095.486p 0.654194mV 82112.02p 0.676494mV 82119.805p 0.672906mV 82124.906p 0.663861mV 82134.227p 0.65428mV 82148.97p 0.597985mV 82160.458p 0.56457mV 82160.747p 0.56457mV 82179.852p 0.5261mV 82180.971p 0.521641mV 82191.791p 0.518545mV 82218.721p 0.408998mV 82227.392p 0.374957mV 83010.048p 0.561179mV 83011.223p 0.561179mV 83022.34p 0.528219mV 83025.437p 0.514911mV 83044.421p 0.448588mV 83066.46p 0.368726mV 84013.686p 0.558719mV 84017.66p 0.558332mV 84040.977p 0.474661mV 84071.173p 0.338656mV 84076.886p 0.332061mV 85009.944p 0.550951mV 85021.363p 0.548957mV 85067.852p 0.504191mV 85086.032p 0.45936mV 87000.016p 0.549333mV 88079.435p 0.511311mV 88106.677p 0.473481mV 88155.329p 0.596284mV 88163.769p 0.64016mV 89000.445p 0.561192mV 89009.138p 0.560166mV 89021.271p 0.519638mV 89027.872p 0.493493mV 89046.367p 0.372643mV 90007.754p 0.596393mV 90018.62p 0.589481mV 90030.188p 0.590454mV 90033.896p 0.590454mV 90054.471p 0.595002mV 90055.11p 0.609332mV 90062.192p 0.61765mV 90088.356p 0.571008mV 90094.255p 0.543872mV 90112.264p 0.485548mV 91077.346p 0.507739mV 91079.158p 0.507739mV 91094.792p 0.581457mV 91120.784p 0.741055mV 92001.963p 0.542293mV 92013.861p 0.548936mV 92015.987p 0.549035mV 93051.393p 0.442555mV 93072.05p 0.398049mV 93076.187p 0.391105mV 94023.079p 0.507502mV 94061.159p 0.397604mV 94108.676p 0.355992mV 94118.621p 0.356228mV 94130.631p 0.36303mV 94131.105p 0.36303mV 94132.293p 0.36303mV 94148.031p 0.365434mV 95007.348p 0.537178mV 95017.23p 0.556974mV 95022.057p 0.563643mV 95041.88p 0.64179mV 95046.757p 0.668389mV 95065.209p 0.756854mV 95065.873p 0.756854mV 96023.009p 0.636211mV 96053.123p 0.725071mV 96070.623p 0.74571mV 96083.722p 0.750673mV 96090.638p 0.760543mV 96092.148p 0.760543mV 97003.07p 0.553197mV 97004.323p 0.553197mV 97007.409p 0.554222mV 97018.103p 0.550038mV 97018.804p 0.550038mV 97025.301p 0.533263mV 97062.631p 0.487199mV 97064.214p 0.487199mV 97079.407p 0.466529mV 97083.234p 0.471237mV 97086.519p 0.481699mV 97111.761p 0.483343mV 97133.052p 0.487296mV 97134.564p 0.487296mV 97160.48p 0.385922mV 97162.377p 0.385922mV 98014.566p 0.53758mV 98030.088p 0.583663mV 98043.709p 0.638615mV 98049.569p 0.663416mV 98060.422p 0.729178mV 98062.249p 0.729178mV 98064.264p 0.729178mV 98068.627p 0.744577mV 98076.652p 0.772613mV 99011.859p 0.511753mV 99012.232p 0.511753mV 99014.294p 0.511753mV 99036.509p 0.637308mV 100023.62p 0.564996mV 100025.092p 0.590391mV 100084.707p 0.762986mV 101000.838p 0.560454mV 101013.678p 0.552793mV 101021.115p 0.545339mV 101066.614p 0.422248mV 101074.065p 0.40046mV 101099.751p 0.358337mV 102007.686p 0.589954mV 102026.114p 0.570553mV 102042.787p 0.551268mV 102059.43p 0.513472mV 102076.833p 0.418445mV 102088.952p 0.386356mV 102090.799p 0.365849mV 103042.371p 0.695967mV 104006.468p 0.507055mV 104017.899p 0.501295mV 104041.224p 0.5545mV 104057.612p 0.569971mV 104061.174p 0.562735mV 104061.507p 0.562735mV 104066.514p 0.549325mV 104067.716p 0.549325mV 104071.34p 0.542296mV 104120.985p 0.538141mV 104137.383p 0.527177mV 104170.884p 0.575474mV 104175.726p 0.585833mV 104189.781p 0.600795mV 104201.728p 0.622176mV 104229.896p 0.611531mV 104250.892p 0.654859mV 104252.733p 0.654859mV 104260.857p 0.694319mV 104266.968p 0.712014mV 104269.524p 0.712014mV 104278.105p 0.743973mV 104288.809p 0.767959mV 104309.185p 0.757868mV 104313.777p 0.755712mV 104357.518p 0.750293mV 104367.13p 0.75439mV 104368.625p 0.75439mV 104373.527p 0.767576mV 105003.655p 0.533546mV 105020.522p 0.532743mV 105039.549p 0.524512mV 105043.62p 0.529901mV 105053.594p 0.559132mV 105054.888p 0.559132mV 105067.352p 0.587114mV 105094.486p 0.57879mV 105111.733p 0.530441mV 105130.209p 0.393073mV 106003.109p 0.565836mV 106023.308p 0.537837mV 106077.281p 0.426077mV 106080.227p 0.403067mV 106081.346p 0.403067mV 107016.633p 0.569129mV 107027.965p 0.525146mV 107054.063p 0.479081mV 107054.76p 0.479081mV 107056.555p 0.477607mV 107096.15p 0.43546mV 107127.074p 0.4428mV 107165.141p 0.528861mV 107171.063p 0.545505mV 107176.193p 0.568317mV 107196.039p 0.673436mV 107199.308p 0.673436mV 107200.24p 0.691434mV 107204.363p 0.691434mV 107211.902p 0.711117mV 108015.98p 0.583548mV 109001.51p 0.51085mV 109009.245p 0.510864mV 109023.827p 0.471605mV 109047.147p 0.334228mV 110037.775p 0.485582mV 110038.143p 0.485582mV 110070.195p 0.457835mV 111000.453p 0.560072mV 111003.77p 0.560072mV 111012.486p 0.555912mV 111029.192p 0.527962mV 111052.375p 0.512742mV 111054.369p 0.512742mV 112029.364p 0.538867mV 112039.98p 0.505971mV 112058.144p 0.411894mV 113002.801p 0.57291mV 113003.085p 0.57291mV 113030.35p 0.59977mV 113039.576p 0.601727mV 113056.308p 0.549686mV 114009.72p 0.514822mV 114041.056p 0.482074mV 114084.684p 0.500056mV 114101.949p 0.510811mV 114110.169p 0.527206mV 114130.329p 0.608642mV 114144.291p 0.650228mV 115035.004p 0.627058mV 115038.868p 0.627058mV 115043.632p 0.623466mV 115053.75p 0.611434mV 115067.755p 0.643642mV 115070.145p 0.667833mV 115083.557p 0.724414mV 115088.664p 0.744638mV 115093.881p 0.772159mV 116018.443p 0.545574mV 116034.293p 0.545446mV 116068.224p 0.653813mV 116096.12p 0.718639mV 116096.226p 0.718639mV 116096.248p 0.718639mV 116112.555p 0.717217mV 116126.272p 0.731412mV 116146.624p 0.765684mV 118030.771p 0.561211mV 118052.361p 0.687069mV 118056.567p 0.725909mV 119014.738p 0.501964mV 119028.64p 0.491197mV 119064.611p 0.467425mV 120012.978p 0.592442mV 120023.671p 0.610906mV 120030.453p 0.61812mV 120033.431p 0.61812mV 120036.868p 0.63174mV 120048.756p 0.679206mV 120052.046p 0.713243mV 120058.426p 0.741833mV 121009.609p 0.542756mV 121023.509p 0.505253mV 121032.126p 0.473202mV 121048.448p 0.412531mV 121053.176p 0.403474mV 121060.434p 0.363995mV 121068.082p 0.345882mV 122024.598p 0.554508mV 122026.905p 0.529593mV 123059.798p 0.358259mV 124039.975p 0.65303mV 124044.813p 0.673068mV 124048.319p 0.687483mV 124056.099p 0.699969mV 125018.048p 0.551344mV 125020.632p 0.53218mV 125056.483p 0.441706mV 125056.951p 0.441706mV 125088.948p 0.354723mV 126014.614p 0.555642mV 126015.294p 0.55547mV 126030.082p 0.54252mV 126033.868p 0.54252mV 126074.841p 0.489892mV 127017.76p 0.580317mV 127021.842p 0.598769mV 128005.465p 0.544421mV 128052.585p 0.73431mV 128057.793p 0.762951mV 129000.917p 0.517191mV 129025.244p 0.51927mV 129028.34p 0.51927mV 129048.881p 0.454004mV 130011.103p 0.585528mV 130013.537p 0.585528mV 130061.507p 0.591879mV 130085.621p 0.533309mV 130087.163p 0.533309mV 130096.86p 0.508889mV 130099.028p 0.508889mV 130100.965p 0.505874mV 130115.413p 0.49515mV 130119.896p 0.49515mV 130127.185p 0.492593mV 131020.693p 0.557526mV 131026.489p 0.570413mV 131033.21p 0.577045mV 131034.692p 0.577045mV 131048.23p 0.597927mV 131060.229p 0.564587mV 131066.886p 0.541359mV 131068.741p 0.541359mV 131087.923p 0.51111mV 131108.155p 0.502654mV 131118.336p 0.47188mV 131136.222p 0.4047mV 132073.243p 0.44161mV 132087.633p 0.421483mV 132088.226p 0.421483mV 132120.609p 0.475332mV 132210.676p 0.555208mV 132217.116p 0.565311mV 133005.715p 0.538753mV 133012.195p 0.544809mV 133023.762p 0.57565mV 133046.325p 0.741287mV 134044.589p 0.480457mV 135036.285p 0.572502mV 135055.902p 0.505833mV 135073.343p 0.423011mV 135080.087p 0.354525mV 136003.103p 0.519609mV 136027.28p 0.476398mV 136051.667p 0.44221mV 136065.158p 0.481732mV 136082.331p 0.547907mV 136095.22p 0.631665mV 137000.832p 0.525507mV 137016.061p 0.52929mV 137020.516p 0.53447mV 137032.941p 0.538171mV 137053.189p 0.557347mV 137100.278p 0.66021mV 138009.987p 0.563676mV 138011.08p 0.569197mV 138017.165p 0.568502mV 138037.441p 0.541572mV 138072.062p 0.472957mV 138096.912p 0.45642mV 138105.47p 0.489375mV 138123.477p 0.519632mV 138193.225p 0.375036mV 139014.252p 0.4903mV 139020.084p 0.495346mV 139043.536p 0.513697mV 139056.401p 0.524554mV 139062.009p 0.527845mV 139092.324p 0.475026mV 139102.0p 0.446985mV 139107.79p 0.429017mV 139116.32p 0.397309mV 140003.892p 0.569723mV 140007.617p 0.569731mV 140010.866p 0.563562mV 141014.254p 0.574678mV 141019.364p 0.588081mV 141034.415p 0.616924mV 141037.943p 0.618793mV 141060.152p 0.628659mV 141081.965p 0.612858mV 141107.163p 0.548926mV 141113.519p 0.550414mV 141151.793p 0.58864mV 141171.527p 0.598353mV 141186.852p 0.608714mV 141203.788p 0.603137mV 141212.676p 0.569842mV 141234.005p 0.441997mV 141248.406p 0.354577mV 142005.195p 0.566267mV 142026.115p 0.592312mV 142058.93p 0.696573mV 142067.57p 0.748683mV 143006.257p 0.512046mV 143028.128p 0.561377mV 143038.91p 0.591904mV 143044.761p 0.610539mV 143061.327p 0.688754mV 143062.815p 0.688754mV 143062.892p 0.688754mV 144003.401p 0.557509mV 144037.797p 0.597766mV 144044.441p 0.603879mV 144057.092p 0.611549mV 144065.088p 0.608011mV 144067.333p 0.608011mV 144106.821p 0.647292mV 144113.232p 0.659216mV 144131.939p 0.739131mV 145009.566p 0.530055mV 145054.816p 0.352241mV 146004.797p 0.500865mV 146009.475p 0.501319mV 146009.54p 0.501319mV 146032.879p 0.517646mV 146043.289p 0.520925mV 146045.413p 0.531696mV 146047.162p 0.531696mV 146070.071p 0.539769mV 147004.43p 0.509391mV 147035.548p 0.516334mV 147041.49p 0.521534mV 147041.722p 0.521534mV 147046.402p 0.532819mV 147071.835p 0.569249mV 147083.506p 0.598189mV 147088.195p 0.62236mV 147100.023p 0.709912mV 147107.579p 0.748808mV 148015.733p 0.587344mV 148028.042p 0.609625mV 148042.227p 0.654977mV 148043.339p 0.654977mV 148061.216p 0.761605mV 149004.167p 0.593045mV 149007.939p 0.592064mV 149020.768p 0.590767mV 149037.425p 0.560446mV 149059.757p 0.475096mV 149063.817p 0.45643mV 150027.391p 0.534214mV 151022.013p 0.471036mV 151064.321p 0.337562mV 152011.098p 0.605556mV 152017.937p 0.606447mV 153033.387p 0.439087mV 154045.625p 0.594875mV 154059.645p 0.605786mV 154060.794p 0.602278mV 154071.597p 0.615174mV 154095.697p 0.638742mV 154103.793p 0.651237mV 155026.274p 0.593492mV 155036.849p 0.600452mV 155053.789p 0.628983mV 155064.089p 0.65219mV 155070.923p 0.690247mV 155073.979p 0.690247mV 155083.429p 0.756323mV 156016.596p 0.585175mV 156018.386p 0.585175mV 156067.917p 0.463857mV 156089.575p 0.392267mV 156092.495p 0.372421mV 157005.352p 0.572793mV 157007.594p 0.572793mV 157025.302p 0.612865mV 157028.55p 0.612865mV 157037.099p 0.65975mV 157039.221p 0.65975mV 158012.681p 0.608554mV 158028.673p 0.667623mV 158035.441p 0.716008mV 158040.19p 0.738318mV 160017.652p 0.564772mV 160018.625p 0.564772mV 160021.358p 0.570721mV 160029.391p 0.583065mV 160032.032p 0.589238mV 160034.78p 0.589238mV 160048.613p 0.621801mV 160060.152p 0.638902mV 160080.065p 0.677756mV 160086.202p 0.68294mV 160105.284p 0.774673mV 161025.753p 0.551831mV 161038.729p 0.557518mV 161062.956p 0.575425mV 161100.243p 0.592755mV 161110.312p 0.58967mV 161166.759p 0.424279mV 161174.06p 0.429019mV 161201.102p 0.498674mV 161214.286p 0.542774mV 161237.258p 0.712371mV 161240.039p 0.763967mV 161244.597p 0.763967mV 162000.3p 0.561261mV 162006.266p 0.560771mV 162014.251p 0.566655mV 162029.892p 0.559616mV 162031.779p 0.553234mV 162032.988p 0.553234mV 163025.46p 0.579643mV 163035.498p 0.573695mV 163076.27p 0.515794mV 164041.921p 0.40979mV 164060.753p 0.337872mV 165001.664p 0.54786mV 165006.966p 0.547002mV 166006.719p 0.595355mV 166013.232p 0.601178mV 166016.29p 0.613581mV 167023.046p 0.598577mV 167025.514p 0.624877mV 167047.411p 0.760211mV 168005.409p 0.539062mV 168008.906p 0.539062mV 168017.98p 0.520128mV 168020.964p 0.501067mV 168039.932p 0.454913mV 168050.267p 0.423143mV 168061.556p 0.396336mV 169020.917p 0.550222mV 169072.24p 0.480223mV 169077.506p 0.478185mV 169082.055p 0.469421mV 169088.309p 0.453918mV 169089.958p 0.453918mV 169108.48p 0.398197mV 170010.694p 0.590263mV 170029.396p 0.583603mV 170046.999p 0.523066mV 170048.655p 0.523066mV 171008.079p 0.522672mV 172022.383p 0.521519mV 172027.656p 0.520346mV 172033.357p 0.512695mV 172048.03p 0.488469mV 172065.363p 0.476661mV 173009.939p 0.534843mV 173011.008p 0.527505mV 173031.271p 0.547333mV 173031.404p 0.547333mV 173074.94p 0.405137mV 174006.552p 0.496728mV 174007.96p 0.496728mV 174015.59p 0.514049mV 174045.991p 0.522363mV 174155.915p 0.402336mV 174172.395p 0.39418mV 174192.775p 0.353106mV 175017.257p 0.500307mV 175040.738p 0.438721mV 175063.629p 0.348536mV 176031.308p 0.616112mV 176041.475p 0.637409mV 176079.078p 0.760267mV 177012.032p 0.495427mV 177030.45p 0.44914mV 177040.158p 0.423198mV 178002.349p 0.498067mV 179003.425p 0.551113mV 180042.668p 0.592792mV 180070.843p 0.64355mV 180073.462p 0.64355mV 180081.045p 0.672518mV 180091.486p 0.67918mV 181013.089p 0.56825mV 181075.316p 0.461493mV 181089.184p 0.474445mV 181125.202p 0.573521mV 182002.849p 0.566903mV 182018.987p 0.584349mV 182035.639p 0.673384mV 182037.99p 0.673384mV 182043.635p 0.693708mV 182051.09p 0.730532mV 182063.105p 0.771357mV 183006.104p 0.573325mV 183014.101p 0.568158mV 183022.579p 0.551934mV 183031.81p 0.548525mV 183035.019p 0.549998mV 183039.847p 0.549998mV 183061.783p 0.576595mV 183067.11p 0.578392mV 183159.574p 0.505654mV 183160.383p 0.483859mV 184015.333p 0.501199mV 184028.967p 0.507067mV 184048.201p 0.528191mV 184079.135p 0.574818mV 184085.418p 0.578254mV 184086.306p 0.578254mV 184130.263p 0.555291mV 184138.472p 0.53068mV 184144.773p 0.512405mV 185030.083p 0.525963mV 185033.598p 0.525963mV 185067.936p 0.441126mV 185068.062p 0.441126mV 186004.263p 0.596007mV 186023.98p 0.596426mV 186028.977p 0.584735mV 186037.931p 0.568447mV 186042.922p 0.551152mV 186067.862p 0.406918mV 186075.88p 0.336752mV 187006.29p 0.515906mV 187010.07p 0.522816mV 187012.15p 0.522816mV 187016.621p 0.535809mV 187019.808p 0.535809mV 187032.436p 0.56145mV 187060.892p 0.710319mV 188054.177p 0.334958mV 189001.213p 0.501211mV 189017.562p 0.508414mV 189021.846p 0.501852mV 189025.881p 0.488733mV 190019.439p 0.590394mV 190036.544p 0.595802mV 190055.478p 0.567519mV 190102.004p 0.578347mV 190111.016p 0.592454mV 190135.066p 0.692578mV 190141.021p 0.717991mV 190146.717p 0.738057mV 191033.393p 0.415132mV 191038.942p 0.386961mV 192002.803p 0.501281mV 192087.58p 0.424573mV 192108.65p 0.394881mV 192112.215p 0.388423mV 193000.172p 0.526538mV 194001.188p 0.576139mV 194004.713p 0.576139mV 194026.752p 0.628897mV 194056.212p 0.754274mV 194063.361p 0.767095mV 195002.378p 0.500322mV 195014.887p 0.507005mV 195025.364p 0.562108mV 195030.14p 0.580176mV 195040.445p 0.597752mV 195085.555p 0.688117mV 195094.171p 0.711804mV 196002.643p 0.524168mV 196026.373p 0.489466mV 197009.789p 0.519312mV 197026.229p 0.490694mV 197034.582p 0.495353mV 197043.53p 0.484703mV 197055.896p 0.431205mV 197094.004p 0.421479mV 197102.109p 0.406932mV 197103.724p 0.406932mV 197111.682p 0.376467mV 198037.487p 0.603982mV 198059.854p 0.606837mV 198069.431p 0.616743mV 198115.733p 0.757748mV 199028.248p 0.500219mV 199047.418p 0.50612mV 199059.404p 0.494799mV 199062.394p 0.49811mV 199106.134p 0.363771mV 199114.813p 0.336358mV 200034.24p 0.5248mV 200042.709p 0.490391mV 200055.177p 0.452323mV 200059.156p 0.452323mV 200067.567p 0.413949mV 200084.745p 0.38502mV 200086.853p 0.365216mV 201021.126p 0.6037mV 201059.739p 0.734268mV 202011.111p 0.539686mV 202035.305p 0.525405mV 202076.222p 0.371539mV 203024.075p 0.605528mV 203027.967p 0.607585mV 203031.581p 0.616285mV 203034.453p 0.616285mV 203038.408p 0.631639mV 203041.508p 0.641122mV 203073.932p 0.754661mV 203074.747p 0.754661mV 204034.864p 0.471943mV 204037.983p 0.445984mV 204038.093p 0.445984mV 204040.128p 0.413253mV 205017.184p 0.512826mV 205025.438p 0.52835mV 205026.972p 0.52835mV 205037.226p 0.543094mV 205079.314p 0.704372mV 205081.011p 0.735931mV 205084.024p 0.735931mV 205088.249p 0.774677mV 205089.215p 0.774677mV 205089.752p 0.774677mV 206023.186p 0.563031mV 206035.422p 0.568563mV 206062.951p 0.499541mV 206069.908p 0.486754mV 206086.436p 0.444329mV 207014.172p 0.588049mV 207017.651p 0.589395mV 207018.287p 0.589395mV 207043.924p 0.631672mV 207045.774p 0.634946mV 207088.163p 0.746405mV 208117.501p 0.691824mV 208131.459p 0.731771mV 208148.344p 0.762749mV 209011.477p 0.582058mV 209017.99p 0.581476mV 209052.576p 0.583745mV 209070.691p 0.564902mV 209080.46p 0.53733mV 210011.295p 0.595793mV 210040.723p 0.578238mV 210045.105p 0.568736mV 210092.768p 0.528048mV 210097.681p 0.530518mV 210116.637p 0.526682mV 210148.147p 0.478693mV 210164.718p 0.452746mV 210182.568p 0.430866mV 210194.027p 0.428044mV 211010.024p 0.525128mV 211014.609p 0.525128mV 211090.114p 0.482561mV 211108.076p 0.496075mV 212040.987p 0.677962mV 212047.863p 0.681587mV 212067.693p 0.729616mV 213005.749p 0.501085mV 213019.795p 0.495612mV 214003.494p 0.51677mV 214004.316p 0.51677mV 214021.394p 0.474964mV 214043.859p 0.326262mV 214044.116p 0.326262mV 215003.441p 0.557631mV 215027.645p 0.533284mV 215035.168p 0.502047mV 215038.161p 0.502047mV 215051.112p 0.475465mV 215067.998p 0.451505mV 215101.483p 0.405275mV 215110.794p 0.394534mV 215135.131p 0.39761mV 215167.005p 0.325008mV 216003.28p 0.508685mV 216012.57p 0.513424mV 216032.605p 0.532544mV 216095.67p 0.675244mV 216107.798p 0.709068mV 216114.819p 0.730391mV 217061.272p 0.48654mV 218013.364p 0.50949mV 218015.272p 0.520629mV 218043.809p 0.592591mV 218060.18p 0.687648mV 218068.99p 0.712757mV 218072.11p 0.744969mV 219001.97p 0.597424mV 219043.267p 0.498569mV 220009.925p 0.520538mV 220010.834p 0.513303mV 220080.601p 0.459503mV 220098.998p 0.492904mV 220127.476p 0.64583mV 220140.829p 0.73586mV 221036.326p 0.559574mV 221044.874p 0.553682mV 221045.918p 0.541548mV 221055.216p 0.510973mV 221087.212p 0.54015mV 221105.809p 0.535427mV 221131.178p 0.508372mV 221146.135p 0.532065mV 221148.369p 0.532065mV 221199.93p 0.530905mV 221200.986p 0.520964mV 222042.923p 0.60759mV 222051.674p 0.606583mV 222080.308p 0.688822mV 222082.323p 0.688822mV 222083.411p 0.688822mV 222091.213p 0.721397mV 222093.644p 0.721397mV 223008.554p 0.497406mV 223046.922p 0.610599mV 223052.644p 0.615655mV 223058.945p 0.614802mV 223063.144p 0.608074mV 223074.853p 0.576933mV 223075.609p 0.55239mV 223077.367p 0.55239mV 223099.213p 0.391193mV 224016.328p 0.505475mV 224034.665p 0.464609mV 225015.739p 0.508795mV 225050.98p 0.433688mV 226023.786p 0.590843mV 226034.237p 0.611963mV 226042.376p 0.634415mV 226069.181p 0.76626mV 227009.916p 0.597629mV 227012.364p 0.591851mV 227100.654p 0.470943mV 228037.679p 0.488919mV 229076.896p 0.4989mV 229134.478p 0.634647mV 230007.381p 0.568695mV 230021.557p 0.569878mV 230055.803p 0.517924mV 230065.049p 0.524288mV 230100.465p 0.595987mV 230172.748p 0.426207mV 230200.727p 0.389294mV 230201.466p 0.389294mV 230203.236p 0.389294mV 231002.862p 0.589674mV 231025.366p 0.60365mV 231035.575p 0.637429mV 231038.404p 0.637429mV 231053.644p 0.694892mV 231054.439p 0.694892mV 231072.678p 0.753796mV 232000.792p 0.527129mV 232026.397p 0.464445mV 232027.916p 0.464445mV 232044.321p 0.385031mV 233000.258p 0.535406mV 233044.023p 0.501127mV 233046.197p 0.486727mV 234017.65p 0.598109mV 234025.96p 0.59223mV 234035.403p 0.574855mV 234047.204p 0.570962mV 234078.466p 0.549472mV 234093.797p 0.555009mV 234106.564p 0.516734mV 234127.018p 0.459483mV 235025.343p 0.507815mV 235042.543p 0.503245mV 236015.158p 0.56596mV 236017.315p 0.56596mV 236019.474p 0.56596mV 236026.641p 0.583819mV 236047.62p 0.596479mV 236056.202p 0.591823mV 236065.426p 0.588238mV 236107.558p 0.609339mV 236136.13p 0.707623mV 236141.396p 0.733463mV 236149.375p 0.766511mV 237036.998p 0.637531mV 237048.658p 0.663292mV 237056.734p 0.679006mV 237065.477p 0.672781mV 237077.698p 0.669754mV 237090.915p 0.636512mV 237113.573p 0.634084mV 237151.949p 0.719004mV 238030.677p 0.505353mV 238037.577p 0.504573mV 238048.348p 0.508461mV 238048.879p 0.508461mV 238094.188p 0.369038mV 239036.563p 0.608925mV 240017.034p 0.558455mV 240026.338p 0.538645mV 240032.662p 0.519324mV 240045.168p 0.473089mV 240059.438p 0.463546mV 240067.013p 0.451911mV 240086.981p 0.446586mV 240087.653p 0.446586mV 241007.125p 0.557262mV 241021.289p 0.555031mV 241060.175p 0.525421mV 242056.285p 0.463549mV 242075.143p 0.424833mV 242154.814p 0.355329mV 243000.666p 0.519999mV 243030.435p 0.496783mV 243032.226p 0.496783mV 243036.281p 0.482581mV 244006.592p 0.597078mV 244029.335p 0.534062mV 244029.599p 0.534062mV 244029.781p 0.534062mV 244031.696p 0.502948mV 244034.058p 0.502948mV 244040.542p 0.459123mV 244096.865p 0.444064mV 244100.083p 0.441546mV 245021.363p 0.601115mV 245031.714p 0.621329mV 245043.66p 0.630538mV 245059.308p 0.657349mV 245074.948p 0.695812mV 245088.009p 0.74804mV 246042.376p 0.659223mV 246058.402p 0.698583mV 246068.829p 0.739334mV 246071.377p 0.751919mV 247021.506p 0.602038mV 247022.003p 0.602038mV 247031.177p 0.611295mV 247048.805p 0.624705mV 247052.524p 0.634213mV 247056.836p 0.650475mV 248002.706p 0.520123mV 248005.002p 0.52047mV 248050.991p 0.403323mV 248051.489p 0.403323mV 248058.462p 0.386882mV 249014.502p 0.585333mV 249052.754p 0.757908mV 250007.967p 0.59024mV 250041.614p 0.57814mV 250049.785p 0.566509mV 250058.361p 0.550002mV 250065.931p 0.533742mV 250075.27p 0.517317mV 250076.651p 0.517317mV 250120.533p 0.432138mV 250150.128p 0.407226mV 250150.241p 0.407226mV 250182.562p 0.386591mV 250218.166p 0.382439mV 250241.603p 0.381313mV 251009.372p 0.49994mV 251044.522p 0.462513mV 251100.988p 0.544118mV 251116.54p 0.579565mV 251149.892p 0.750057mV 252059.183p 0.566729mV 252060.035p 0.573279mV 252077.378p 0.606368mV 252078.206p 0.606368mV 252097.376p 0.688654mV 252118.065p 0.770095mV 253002.997p 0.540775mV 253007.055p 0.540161mV 253013.758p 0.54579mV 253023.893p 0.575803mV 253037.57p 0.59314mV 253040.148p 0.586811mV 253050.104p 0.568636mV 253056.351p 0.569268mV 253063.943p 0.563716mV 253077.977p 0.509804mV 253083.772p 0.479168mV 253104.511p 0.377433mV 254028.503p 0.549341mV 254040.365p 0.55984mV 254041.38p 0.55984mV 254043.281p 0.55984mV 254062.392p 0.544931mV 254112.08p 0.702194mV 254116.838p 0.729734mV 255029.709p 0.596896mV 255035.828p 0.61962mV 255066.947p 0.698716mV 255075.802p 0.730828mV 255080.614p 0.745253mV 256047.097p 0.601583mV 256068.751p 0.650697mV 256117.549p 0.675067mV 256142.878p 0.69037mV 256158.813p 0.642703mV 256170.47p 0.557474mV 256178.551p 0.525543mV 257027.533p 0.536213mV 257029.379p 0.536213mV 257055.705p 0.430267mV 257062.369p 0.410093mV 257063.345p 0.410093mV 258035.663p 0.659243mV 258036.533p 0.659243mV 258046.035p 0.696332mV 258055.008p 0.711665mV 258062.48p 0.723881mV 259053.931p 0.527364mV 259071.882p 0.540102mV 259128.532p 0.556583mV 259159.182p 0.501644mV 259184.087p 0.41841mV 260007.654p 0.526284mV 261039.323p 0.589552mV 261084.227p 0.672242mV 262090.382p 0.623215mV 262091.857p 0.623215mV 262094.1p 0.623215mV 262100.351p 0.677151mV 262108.005p 0.701823mV 263005.688p 0.559715mV 263017.901p 0.542343mV 263048.192p 0.540077mV 263079.209p 0.548121mV 263116.307p 0.434684mV 264025.672p 0.625221mV 264079.908p 0.617102mV 264104.921p 0.554201mV 264124.903p 0.541152mV 264129.19p 0.525319mV 264137.468p 0.512289mV 264140.277p 0.514928mV 264167.616p 0.518761mV 265014.216p 0.51694mV 265032.584p 0.54233mV 265038.879p 0.554612mV 265052.059p 0.616724mV 265093.842p 0.763708mV 265096.591p 0.771151mV 266034.8p 0.412101mV 266043.319p 0.386114mV 266054.869p 0.356314mV 267030.089p 0.588957mV 267035.962p 0.61378mV 267035.993p 0.61378mV 267048.591p 0.645432mV 267067.016p 0.71566mV 268003.423p 0.577187mV 268026.722p 0.594152mV 268044.411p 0.599716mV 268045.982p 0.60222mV 268054.021p 0.598744mV 268058.808p 0.60189mV 268061.067p 0.599049mV 268073.683p 0.588039mV 268086.286p 0.582861mV 268090.861p 0.594115mV 268106.155p 0.629356mV 268118.598p 0.648442mV 268127.919p 0.644698mV 268131.853p 0.634355mV 268146.966p 0.606667mV 268147.549p 0.606667mV 268149.255p 0.606667mV 268175.814p 0.593214mV 268183.035p 0.599267mV 268208.264p 0.666144mV 268214.702p 0.687321mV 269038.005p 0.528428mV 269049.441p 0.532954mV 269052.128p 0.538198mV 269053.095p 0.538198mV 269068.446p 0.540777mV 269079.295p 0.519074mV 269079.468p 0.519074mV 269083.11p 0.498635mV 270025.575p 0.5829mV 270041.764p 0.648769mV 270054.812p 0.696965mV 270058.322p 0.725275mV 270063.755p 0.748267mV 271001.898p 0.586966mV 271002.489p 0.586966mV 271013.273p 0.591416mV 271038.947p 0.629476mV 271047.685p 0.651223mV 272011.125p 0.539829mV 272045.492p 0.5187mV 272049.41p 0.5187mV 272064.513p 0.515506mV 272068.241p 0.501498mV 272077.103p 0.453852mV 272120.555p 0.355792mV 273000.512p 0.58032mV 273017.671p 0.577559mV 273058.909p 0.529339mV 273064.603p 0.512252mV 273073.484p 0.471278mV 273073.763p 0.471278mV 273080.21p 0.441395mV 273091.611p 0.409207mV 274038.291p 0.617589mV 275005.613p 0.56823mV 275015.156p 0.574959mV 275018.966p 0.574959mV 275029.651p 0.59487mV 275057.157p 0.688603mV 275062.008p 0.686849mV 275088.434p 0.697065mV 275090.975p 0.700403mV 275091.586p 0.700403mV 275100.835p 0.728573mV 275104.572p 0.728573mV 276007.326p 0.599865mV 276033.368p 0.585093mV 276052.947p 0.629984mV 276053.781p 0.629984mV 277022.982p 0.552277mV 277051.232p 0.494545mV 277070.49p 0.4503mV 278006.567p 0.554966mV 278030.722p 0.637369mV 278051.273p 0.707895mV 279009.284p 0.548034mV 279016.456p 0.552594mV 279029.998p 0.557202mV 279058.189p 0.444551mV 280009.626p 0.549999mV 280028.899p 0.500543mV 280054.802p 0.464297mV 280075.256p 0.484381mV 280099.24p 0.575685mV 280102.397p 0.601198mV 280123.712p 0.731717mV 281009.733p 0.571402mV 281013.568p 0.564667mV 281030.96p 0.538538mV 281031.521p 0.538538mV 281050.603p 0.498986mV 281050.805p 0.498986mV 281074.832p 0.493224mV 281075.694p 0.49101mV 281077.166p 0.49101mV 281152.386p 0.42746mV 281157.432p 0.425345mV 281171.419p 0.439372mV 281195.19p 0.381179mV 282004.071p 0.516507mV 282012.511p 0.509421mV 282016.679p 0.496112mV 282020.721p 0.476251mV 282023.879p 0.476251mV 282029.647p 0.462344mV 282033.239p 0.454258mV 282036.249p 0.451898mV 282063.088p 0.399549mV 283011.071p 0.568105mV 283013.872p 0.568105mV 283018.67p 0.567473mV 283056.761p 0.670147mV 283067.196p 0.718936mV 283067.357p 0.718936mV 283070.658p 0.753955mV 283071.043p 0.753955mV 284036.352p 0.567883mV 284044.648p 0.585933mV 284069.062p 0.686227mV 285010.95p 0.594568mV 285016.821p 0.594762mV 285025.178p 0.589699mV 285043.904p 0.606098mV 285056.532p 0.656875mV 285092.354p 0.732731mV 286010.134p 0.596276mV 286048.84p 0.572846mV 286050.399p 0.568574mV 286053.376p 0.568574mV 286079.807p 0.516832mV 287010.31p 0.548424mV 287011.371p 0.548424mV 288016.264p 0.513743mV 288019.985p 0.513743mV 288045.474p 0.507073mV 288045.802p 0.507073mV 288097.299p 0.707497mV 288105.614p 0.750562mV 288105.673p 0.750562mV 289030.555p 0.509758mV 289055.35p 0.501468mV 289075.456p 0.527791mV 289091.961p 0.54224mV 289097.1p 0.551064mV 289118.049p 0.535815mV 289136.567p 0.545117mV 289145.632p 0.530674mV 289214.443p 0.419778mV 289219.24p 0.410239mV 290011.848p 0.536958mV 290033.263p 0.512138mV 290084.491p 0.326475mV 291009.506p 0.592356mV 291017.33p 0.573271mV 292002.296p 0.553216mV 292005.447p 0.552843mV 292033.745p 0.494009mV 292044.008p 0.447867mV 293005.211p 0.533617mV 293007.228p 0.533617mV 294001.6p 0.587283mV 294006.235p 0.586575mV 294023.48p 0.623668mV 294031.064p 0.656351mV 295022.503p 0.547013mV 295023.271p 0.547013mV 295040.997p 0.582575mV 295041.986p 0.582575mV 295063.71p 0.721124mV 296010.611p 0.494889mV 296080.302p 0.348391mV 297008.46p 0.603196mV 298030.668p 0.547589mV 298040.699p 0.555979mV 298041.49p 0.555979mV 298059.198p 0.540278mV 298069.807p 0.523555mV 298102.219p 0.462777mV 298155.885p 0.394044mV 298194.388p 0.366909mV 298200.965p 0.374946mV 298210.398p 0.378547mV 298211.333p 0.378547mV 298245.098p 0.474115mV 298252.233p 0.489877mV 298276.189p 0.633239mV 298279.396p 0.633239mV 298302.499p 0.766052mV 298302.714p 0.766052mV 299053.167p 0.508555mV 299064.813p 0.474026mV 299076.654p 0.422414mV 299079.482p 0.422414mV 299086.949p 0.370128mV 300047.974p 0.637857mV 300051.498p 0.645516mV 301047.175p 0.637242mV 301071.847p 0.762403mV 302002.273p 0.563297mV 302009.141p 0.562403mV 302011.696p 0.567895mV 302049.085p 0.649997mV 303007.908p 0.509737mV 303013.902p 0.516716mV 303040.786p 0.562011mV 303051.25p 0.54393mV 303055.078p 0.544378mV 303073.318p 0.520258mV 304000.477p 0.550135mV 304018.605p 0.572061mV 304029.608p 0.61844mV 305049.449p 0.415445mV 305054.135p 0.392919mV 306009.323p 0.523675mV 306041.717p 0.523872mV 306064.407p 0.586754mV 306086.443p 0.636823mV 306090.212p 0.654253mV 306100.491p 0.672033mV 306101.142p 0.672033mV 306107.875p 0.672587mV 306111.506p 0.667652mV 307032.85p 0.501867mV 307062.732p 0.508006mV 307065.261p 0.504877mV 307077.464p 0.478918mV 308004.963p 0.538537mV 309059.837p 0.482434mV 309077.79p 0.499803mV 309106.472p 0.477647mV 309145.497p 0.576871mV 309150.282p 0.585456mV 309155.146p 0.60051mV 309176.866p 0.651186mV 309179.509p 0.651186mV 309190.614p 0.704172mV 310039.579p 0.508453mV 310076.118p 0.389836mV 310100.457p 0.328174mV 311011.444p 0.5984mV 311016.119p 0.611939mV 312024.84p 0.599228mV 312036.334p 0.645903mV 312074.247p 0.699813mV 312075.198p 0.694978mV 312099.693p 0.659698mV 312102.772p 0.640422mV 312104.482p 0.640422mV 312117.86p 0.561144mV 312123.027p 0.531201mV 312138.59p 0.428409mV 313003.131p 0.601164mV 313046.883p 0.507751mV 313095.413p 0.495477mV 313104.817p 0.498968mV 313107.252p 0.508407mV 313121.113p 0.560247mV 313152.774p 0.621537mV 313152.844p 0.621537mV 313160.189p 0.623821mV 313175.072p 0.614904mV 313209.873p 0.652299mV 313215.74p 0.702146mV 313227.502p 0.76767mV 314006.482p 0.584814mV 314023.09p 0.61434mV 314036.842p 0.640609mV 314040.133p 0.662824mV 314049.497p 0.679331mV 314058.068p 0.720845mV 314062.166p 0.746067mV 314068.039p 0.766143mV 315044.92p 0.394049mV 315046.471p 0.38928mV 315084.567p 0.440859mV 315086.239p 0.441205mV 315109.995p 0.498587mV 315110.127p 0.527234mV 315142.74p 0.717669mV 315143.618p 0.717669mV 316002.05p 0.601481mV 316004.109p 0.601481mV 316005.037p 0.600486mV 316006.613p 0.600486mV 316026.202p 0.574403mV 316052.52p 0.545678mV 316058.037p 0.546128mV 316058.151p 0.546128mV 316060.837p 0.540248mV 316066.174p 0.528042mV 316074.544p 0.509474mV 316090.01p 0.445375mV 317011.486p 0.54448mV 317013.581p 0.54448mV 317014.636p 0.54448mV 317016.503p 0.556081mV 317034.844p 0.55312mV 317048.803p 0.569495mV 317056.632p 0.612171mV 317070.108p 0.71308mV 317072.674p 0.71308mV 318040.289p 0.742895mV 319007.408p 0.581439mV 319057.211p 0.594271mV 319075.785p 0.542906mV 319084.849p 0.514753mV 320003.516p 0.556702mV 320003.592p 0.556702mV 320015.998p 0.563209mV 320032.583p 0.538796mV 321006.018p 0.520125mV 321020.408p 0.509524mV 321073.464p 0.703029mV 321074.583p 0.703029mV 321077.482p 0.729733mV 322001.62p 0.594451mV 322008.416p 0.594735mV 322030.65p 0.644758mV 322031.472p 0.644758mV 322034.998p 0.644758mV 323007.551p 0.530669mV 323011.812p 0.537535mV 323023.107p 0.569846mV 323033.543p 0.589609mV 323038.671p 0.602907mV 323047.827p 0.649223mV 323049.281p 0.649223mV 324021.112p 0.570994mV 324066.884p 0.611336mV 324112.055p 0.671841mV 324135.527p 0.745541mV 325076.737p 0.599634mV 325082.384p 0.598892mV 325101.164p 0.624404mV 325102.02p 0.624404mV 325109.554p 0.63181mV 325111.445p 0.633401mV 325117.725p 0.641788mV 325131.124p 0.670374mV 325142.587p 0.661621mV 325182.771p 0.575323mV 325198.931p 0.604485mV 325206.665p 0.656583mV 325214.432p 0.680148mV 325224.681p 0.748206mV 326025.165p 0.570076mV 326036.664p 0.578911mV 326060.304p 0.60706mV 326077.123p 0.65988mV 326083.95p 0.68268mV 327032.934p 0.572376mV 327060.061p 0.597796mV 327091.945p 0.468337mV 328009.178p 0.571116mV 328098.976p 0.420874mV 329064.896p 0.484765mV 329077.755p 0.451135mV 329087.01p 0.457338mV 329102.836p 0.484124mV 329103.607p 0.484124mV 329115.662p 0.51299mV 329135.472p 0.560564mV 329154.279p 0.630534mV 330004.159p 0.553708mV 330028.029p 0.60271mV 330030.576p 0.609146mV 330033.619p 0.609146mV 330049.248p 0.643232mV 330075.044p 0.696648mV 330079.504p 0.696648mV 330086.809p 0.717078mV 330096.369p 0.716581mV 330108.676p 0.707878mV 330130.866p 0.713178mV 330147.33p 0.676378mV 330153.675p 0.653545mV 330163.038p 0.616346mV 330178.7p 0.51714mV 330181.799p 0.484419mV 331028.9p 0.55265mV 331055.073p 0.666851mV 332020.199p 0.512575mV 332037.19p 0.538933mV 332066.404p 0.57126mV 332107.658p 0.575571mV 332116.285p 0.568756mV 332139.544p 0.632434mV 333002.627p 0.551872mV 333029.102p 0.497213mV 334008.473p 0.567254mV 334052.655p 0.564605mV 334063.423p 0.551177mV 334119.523p 0.363245mV 336020.594p 0.606929mV 336045.133p 0.731984mV 337023.895p 0.524914mV 337063.338p 0.549104mV 337064.487p 0.549104mV 337108.945p 0.58438mV 337112.322p 0.577932mV 337128.608p 0.559693mV 337155.372p 0.620392mV 337174.615p 0.626093mV 337181.239p 0.638613mV 337184.17p 0.638613mV 337196.461p 0.670711mV 337206.213p 0.714139mV 337207.989p 0.714139mV 337252.971p 0.754534mV 337273.679p 0.76112mV 338018.779p 0.546786mV 338037.982p 0.558017mV 338049.114p 0.58867mV 338070.431p 0.596454mV 338073.848p 0.596454mV 338094.798p 0.615155mV 338102.183p 0.61402mV 338135.392p 0.675855mV 338166.997p 0.771493mV 338168.945p 0.771493mV 339020.021p 0.496507mV 339029.634p 0.495074mV 339045.531p 0.43533mV 339046.279p 0.43533mV 339049.344p 0.43533mV 339075.623p 0.345034mV 340045.826p 0.60848mV 340050.921p 0.639711mV 340062.73p 0.722317mV 340069.61p 0.774075mV 341003.307p 0.569556mV 341044.112p 0.503255mV 342013.636p 0.496091mV 342023.61p 0.462084mV 342036.377p 0.398144mV 343000.86p 0.582346mV 343009.383p 0.581319mV 343012.473p 0.574199mV 343036.251p 0.623167mV 343061.026p 0.649896mV 343093.851p 0.609845mV 343096.112p 0.603909mV 343112.959p 0.626009mV 343135.53p 0.77334mV 343137.357p 0.77334mV 344029.114p 0.569886mV 344042.595p 0.587353mV 344057.053p 0.600266mV 344070.494p 0.571681mV 344104.108p 0.460685mV 344110.652p 0.408752mV 345018.403p 0.492448mV 345025.008p 0.51061mV 346003.266p 0.596769mV 346006.246p 0.596769mV 346030.742p 0.556871mV 346031.129p 0.556871mV 346032.775p 0.556871mV 346091.647p 0.363402mV 346108.717p 0.325144mV 347004.531p 0.514834mV 347028.94p 0.51414mV 347032.913p 0.519582mV 347053.073p 0.55214mV 347058.031p 0.550637mV 348038.196p 0.537502mV 348068.204p 0.447931mV 348069.055p 0.447931mV 348097.065p 0.428496mV 349015.496p 0.513832mV 349035.716p 0.410043mV 349040.339p 0.376506mV 349054.324p 0.325304mV 350087.913p 0.402583mV 350096.213p 0.360019mV 350098.182p 0.360019mV 351034.715p 0.570134mV 351036.79p 0.547209mV 352003.985p 0.534143mV 352043.304p 0.498954mV 352047.728p 0.496608mV 352066.098p 0.458564mV 352112.586p 0.449543mV 352116.957p 0.45085mV 352153.228p 0.583234mV 352161.087p 0.623855mV 352163.092p 0.623855mV 353009.47p 0.505181mV 353035.215p 0.43698mV 353038.302p 0.43698mV 353038.533p 0.43698mV 353118.954p 0.391171mV 353120.576p 0.391201mV 353145.292p 0.369801mV 354006.984p 0.504709mV 354023.119p 0.489327mV 354042.973p 0.480706mV 354056.514p 0.488932mV 354102.596p 0.612613mV 354120.993p 0.697169mV 354122.094p 0.697169mV 354123.511p 0.697169mV 355002.179p 0.600962mV 355036.817p 0.610183mV 355046.69p 0.583447mV 355050.055p 0.579984mV 355074.547p 0.593341mV 355095.29p 0.666904mV 355113.024p 0.67575mV 355159.963p 0.68076mV 355161.556p 0.702323mV 356011.81p 0.516085mV 356029.328p 0.522106mV 356046.376p 0.519236mV 356096.37p 0.331108mV 357013.59p 0.509222mV 357013.981p 0.509222mV 357037.024p 0.55582mV 357052.737p 0.590225mV 357062.966p 0.62037mV 357063.304p 0.62037mV 357068.694p 0.645338mV 358030.393p 0.574782mV 358044.874p 0.630778mV 359066.025p 0.674583mV 359071.244p 0.707618mV 359071.5p 0.707618mV 360027.196p 0.456492mV 360044.554p 0.371671mV 361010.178p 0.542096mV 361014.129p 0.542096mV 361014.836p 0.542096mV 361019.244p 0.553541mV 361023.549p 0.558635mV 361028.26p 0.570053mV 361061.0p 0.721068mV 362032.566p 0.635309mV 362035.234p 0.662814mV 362036.393p 0.662814mV 362057.456p 0.754536mV 363010.685p 0.570653mV 363014.904p 0.570653mV 363068.041p 0.516091mV 363070.625p 0.522314mV 363094.194p 0.520063mV 363133.041p 0.58316mV 363140.237p 0.624174mV 363145.385p 0.6357mV 363150.719p 0.641409mV 363155.974p 0.641379mV 363174.777p 0.607047mV 363214.898p 0.411863mV 364006.628p 0.590211mV 364014.037p 0.583573mV 364017.494p 0.570891mV 364063.976p 0.628656mV 365049.438p 0.576826mV 365057.009p 0.582289mV 365082.23p 0.628292mV 365109.849p 0.666016mV 365118.263p 0.694309mV 365126.964p 0.750823mV 366082.762p 0.533564mV 366102.096p 0.635597mV 366110.221p 0.713137mV 367044.283p 0.464052mV 367129.35p 0.616398mV 367153.683p 0.765874mV 368006.061p 0.539819mV 368046.148p 0.49458mV 368046.427p 0.49458mV 368139.783p 0.408402mV 368141.624p 0.404336mV 368148.369p 0.393141mV 369000.317p 0.582632mV 369034.655p 0.615494mV 370011.591p 0.516749mV 370072.134p 0.532586mV 370087.318p 0.612244mV 370093.52p 0.638959mV 371024.145p 0.504087mV 372005.784p 0.497096mV 372009.365p 0.497096mV 372031.073p 0.506043mV 372044.158p 0.518581mV 373001.04p 0.540759mV 373035.924p 0.56571mV 373052.656p 0.58905mV 373079.484p 0.666561mV 373080.398p 0.687328mV 373080.519p 0.687328mV 374021.854p 0.626932mV 374031.514p 0.649962mV 374053.872p 0.703403mV 374083.785p 0.737342mV 374100.65p 0.671806mV 374113.12p 0.650951mV 374134.724p 0.579425mV 374139.59p 0.550044mV 374143.342p 0.527145mV 374147.88p 0.497945mV 374158.459p 0.44524mV 375013.008p 0.570915mV 375015.906p 0.571349mV 375026.132p 0.553713mV 375071.693p 0.439377mV 376035.324p 0.585656mV 376037.352p 0.585656mV 376057.542p 0.61073mV 376099.073p 0.694372mV 376105.161p 0.750477mV 377042.76p 0.450649mV 377134.225p 0.692903mV 378028.845p 0.505997mV 378037.183p 0.483383mV 378057.011p 0.433206mV 378096.614p 0.448187mV 378135.412p 0.456486mV 378190.914p 0.558513mV 378198.503p 0.575913mV 378239.521p 0.75254mV 379074.569p 0.416849mV 379104.254p 0.431947mV 379116.368p 0.419592mV 380011.127p 0.603594mV 380018.113p 0.604753mV 380027.912p 0.614386mV 380031.698p 0.610334mV 380061.256p 0.561324mV 380066.799p 0.552694mV 380097.354p 0.570904mV 380119.276p 0.538207mV 380138.738p 0.492617mV 380149.863p 0.455737mV 380152.592p 0.439801mV 380202.957p 0.469884mV 380240.989p 0.631121mV 380263.021p 0.623439mV 380271.63p 0.610205mV 380273.312p 0.610205mV 380301.034p 0.580093mV 380311.397p 0.559924mV 381055.976p 0.371351mV 381065.742p 0.350805mV 381066.944p 0.350805mV 383021.809p 0.520184mV 383025.969p 0.531874mV 383046.439p 0.5902mV 383076.95p 0.773626mV 384009.004p 0.550635mV 384059.581p 0.755293mV 385002.912p 0.570008mV 385031.181p 0.489348mV 386035.346p 0.510422mV 386061.119p 0.494102mV 386080.994p 0.555673mV 386088.06p 0.576926mV 386102.144p 0.603595mV 386102.471p 0.603595mV 386124.578p 0.592915mV 386129.402p 0.590929mV 387025.38p 0.563381mV 387026.934p 0.563381mV 387031.253p 0.569207mV 387043.997p 0.60005mV 387051.952p 0.644327mV 388001.149p 0.561226mV 388027.975p 0.569575mV 388091.448p 0.706593mV 388154.562p 0.738561mV 388158.85p 0.755732mV 390021.961p 0.556651mV 391023.853p 0.580559mV 391025.384p 0.593762mV 391027.006p 0.593762mV 391031.873p 0.600859mV 391045.111p 0.649207mV 391078.06p 0.756618mV 392024.315p 0.516916mV 392076.886p 0.329483mV 393002.055p 0.589562mV 393012.744p 0.583575mV 393029.278p 0.541645mV 394003.231p 0.502154mV 394003.994p 0.502154mV 394004.411p 0.502154mV 394024.175p 0.498268mV 394101.914p 0.327699mV 395038.196p 0.436713mV 395044.676p 0.415354mV 396043.686p 0.638987mV 396045.124p 0.642041mV 396065.552p 0.697919mV 397013.519p 0.51329mV 397043.737p 0.479852mV 397072.118p 0.330248mV 398002.648p 0.541229mV 398030.263p 0.605323mV 398036.39p 0.617414mV 398037.645p 0.617414mV 398049.681p 0.623847mV 398058.505p 0.606955mV 398076.774p 0.615649mV 398094.583p 0.663924mV 398095.86p 0.681048mV 398137.879p 0.75365mV 399005.984p 0.541327mV 399006.052p 0.541327mV 399027.157p 0.527338mV 399033.071p 0.507989mV 400033.364p 0.623188mV 400048.17p 0.614325mV 400078.828p 0.5753mV 400097.056p 0.537044mV 400131.91p 0.373333mV 400136.131p 0.350739mV 401008.309p 0.528484mV 401023.491p 0.517251mV 401092.921p 0.405161mV 401115.225p 0.434946mV 401119.263p 0.434946mV 401139.162p 0.434782mV 402005.601p 0.574028mV 402010.693p 0.568646mV 402014.505p 0.568646mV 402025.936p 0.55331mV 402042.399p 0.557556mV 402068.857p 0.615807mV 402070.542p 0.62426mV 402088.745p 0.614566mV 402102.703p 0.627776mV 402130.692p 0.64856mV 402165.585p 0.640886mV 402180.576p 0.681564mV 403028.285p 0.554664mV 403095.008p 0.56815mV 403101.29p 0.586mV 403106.297p 0.597663mV 403116.812p 0.602854mV 403118.725p 0.602854mV 403135.566p 0.604711mV 403147.894p 0.601468mV 403151.201p 0.609773mV 403155.647p 0.624696mV 403168.59p 0.649467mV 403192.624p 0.70656mV 403194.735p 0.70656mV 403205.829p 0.738711mV 404026.204p 0.637979mV 405004.301p 0.556218mV 405012.524p 0.564366mV 405015.143p 0.577957mV 405032.147p 0.581777mV 406002.808p 0.587847mV 406009.627p 0.587422mV 406010.892p 0.593533mV 406016.185p 0.606177mV 406030.854p 0.633443mV 406045.063p 0.683805mV 406052.226p 0.693573mV 406077.333p 0.674626mV 406104.693p 0.632893mV 406161.008p 0.478254mV 406168.298p 0.46759mV 406176.696p 0.463691mV 407003.22p 0.49883mV 407012.545p 0.503362mV 407014.989p 0.503362mV 407037.986p 0.557316mV 407083.694p 0.681462mV 407095.879p 0.721135mV 407105.719p 0.750273mV 407106.207p 0.750273mV 407109.95p 0.750273mV 407114.395p 0.763422mV 408001.923p 0.511738mV 408042.747p 0.546514mV 408064.617p 0.5683mV 408084.181p 0.591311mV 408114.621p 0.575881mV 408125.124p 0.574047mV 408145.201p 0.518994mV 408168.238p 0.475347mV 408169.349p 0.475347mV 409028.937p 0.644797mV 409030.799p 0.678227mV 409041.084p 0.765861mV 410007.87p 0.594677mV 411013.31p 0.602773mV 411017.795p 0.616139mV 411057.279p 0.740862mV 411057.377p 0.740862mV 412006.383p 0.51024mV 413031.993p 0.472346mV 413050.524p 0.519182mV 413064.015p 0.54066mV 413087.232p 0.514046mV 413090.932p 0.489653mV 413109.056p 0.439736mV 413115.977p 0.418343mV 413130.677p 0.427281mV 413218.732p 0.640136mV 413225.273p 0.683101mV 414008.718p 0.600856mV 414023.782p 0.629842mV 414032.565p 0.62823mV 414071.685p 0.589931mV 414097.376p 0.522492mV 414144.027p 0.425979mV 414154.874p 0.423699mV 414160.465p 0.405803mV 414180.503p 0.397005mV 414187.245p 0.380084mV 414191.301p 0.355977mV 415037.5p 0.418633mV 416000.435p 0.598987mV 416010.264p 0.604156mV 416017.603p 0.616641mV 416028.952p 0.636417mV 416054.035p 0.730744mV 416059.363p 0.736132mV 416067.473p 0.731743mV 416076.532p 0.744388mV 417022.174p 0.608328mV 417048.078p 0.687031mV 418000.297p 0.504033mV 418014.772p 0.497189mV 418021.444p 0.489144mV 418025.775p 0.487763mV 419003.304p 0.560039mV 419016.469p 0.569124mV 419022.319p 0.576534mV 419030.08p 0.585461mV 419042.617p 0.620324mV 419049.067p 0.647623mV 419052.276p 0.681647mV 419059.77p 0.710008mV 420029.493p 0.570883mV 420049.734p 0.584822mV 420068.545p 0.551373mV 420069.03p 0.551373mV 420102.143p 0.484151mV 421030.2p 0.629913mV 421044.899p 0.64071mV 421075.612p 0.720902mV 421086.092p 0.733249mV 421099.468p 0.762416mV 422006.199p 0.534461mV 422032.946p 0.513944mV 423004.113p 0.5033mV 423006.989p 0.50406mV 423014.815p 0.498231mV 423025.853p 0.466231mV 423091.403p 0.486861mV 423103.472p 0.511697mV 423104.126p 0.511697mV 423130.148p 0.51715mV 423139.062p 0.518469mV 423140.115p 0.525878mV 424021.005p 0.62672mV 424023.175p 0.62672mV 424023.83p 0.62672mV 425008.847p 0.544305mV 425019.414p 0.526271mV 425024.399p 0.50771mV 425030.803p 0.463723mV 425041.321p 0.443232mV 425054.575p 0.445363mV 425055.552p 0.454807mV 425063.173p 0.469861mV 425089.727p 0.557242mV 425105.158p 0.547518mV 425113.659p 0.548304mV 425129.615p 0.550629mV 425165.913p 0.686431mV 425179.829p 0.737402mV 426003.037p 0.574467mV 426028.913p 0.626134mV 426035.715p 0.635109mV 426041.386p 0.63094mV 426086.119p 0.681658mV 426092.929p 0.706895mV 427033.883p 0.584782mV 427036.86p 0.610316mV 427045.023p 0.655894mV 427049.459p 0.655894mV 427061.436p 0.725314mV 428053.275p 0.518848mV 428092.182p 0.644759mV 428110.359p 0.72273mV 428111.316p 0.72273mV 430000.923p 0.562996mV 430049.95p 0.770185mV 431026.191p 0.569391mV 431050.298p 0.532056mV 431075.891p 0.43713mV 432000.708p 0.589533mV 432004.564p 0.589533mV 432010.699p 0.596579mV 432014.392p 0.596579mV 432027.994p 0.618601mV 432039.26p 0.628714mV 432040.417p 0.637609mV 432041.549p 0.637609mV 432067.552p 0.735161mV 432071.099p 0.760992mV 433001.877p 0.49629mV 433003.227p 0.49629mV 433008.447p 0.496271mV 433014.989p 0.48962mV 433032.599p 0.459071mV 433057.519p 0.389854mV 433057.876p 0.389854mV 433063.995p 0.377502mV 433078.603p 0.346598mV 434001.341p 0.52199mV 434008.812p 0.521355mV 434017.887p 0.500653mV 434018.643p 0.500653mV 434022.903p 0.480539mV 434026.338p 0.45382mV 435066.868p 0.331806mV 436015.016p 0.523863mV 436049.073p 0.483726mV 436089.613p 0.499872mV 436108.866p 0.61058mV 436124.824p 0.729789mV 436127.503p 0.762607mV 437007.803p 0.570145mV 437021.445p 0.573334mV 437036.112p 0.521205mV 437076.465p 0.345454mV 438009.724p 0.500254mV 438062.234p 0.478972mV 438102.916p 0.357036mV 439002.911p 0.540567mV 439005.521p 0.540271mV 439006.289p 0.540271mV 439030.862p 0.543958mV 439037.241p 0.555792mV 439081.361p 0.608392mV 439090.336p 0.616042mV 439114.213p 0.636127mV 439166.58p 0.500536mV 440004.31p 0.526893mV 440005.361p 0.525944mV 440040.389p 0.476619mV 440045.714p 0.461438mV 441029.343p 0.548975mV 441032.698p 0.567662mV 441033.734p 0.567662mV 441074.045p 0.764962mV 442055.35p 0.710692mV 443001.075p 0.603414mV 443011.744p 0.598705mV 443016.575p 0.600006mV 443033.566p 0.605747mV 443041.329p 0.604821mV 443063.764p 0.569261mV 443119.974p 0.383215mV 444026.233p 0.502676mV 444028.778p 0.502676mV 444071.119p 0.613811mV 444100.584p 0.642048mV 444101.907p 0.642048mV 444102.388p 0.642048mV 444127.262p 0.606003mV 444138.737p 0.565928mV 445009.674p 0.567201mV 445022.983p 0.55548mV 445046.59p 0.468973mV 447000.267p 0.573057mV 447005.802p 0.573859mV 447013.912p 0.581108mV 447034.336p 0.675236mV 447038.918p 0.702998mV 447047.381p 0.742306mV 448001.327p 0.549843mV 448004.377p 0.549843mV 448029.535p 0.496141mV 448055.256p 0.350244mV 449014.107p 0.593796mV 449018.465p 0.593644mV 449021.553p 0.600064mV 449022.661p 0.600064mV 449025.499p 0.600464mV 449039.042p 0.608506mV 449047.103p 0.592792mV 449063.328p 0.574718mV 449069.701p 0.564925mV 449071.759p 0.548987mV 449118.178p 0.438713mV 449121.641p 0.431265mV 449147.655p 0.350992mV 450004.939p 0.587779mV 451002.153p 0.54977mV 451035.474p 0.527099mV 451038.713p 0.527099mV 451053.476p 0.485694mV 451069.907p 0.384922mV 452009.629p 0.516712mV 452023.872p 0.502368mV 452032.057p 0.506209mV 452070.207p 0.549603mV 452082.485p 0.575381mV 452112.329p 0.669069mV 453001.492p 0.593265mV 453062.566p 0.531333mV 453115.163p 0.554151mV 453118.374p 0.554151mV 453127.341p 0.564481mV 453136.275p 0.562483mV 453138.339p 0.562483mV 453170.196p 0.43917mV 453172.569p 0.43917mV 454000.626p 0.547647mV 454003.57p 0.547647mV 454023.009p 0.510974mV 454048.996p 0.356229mV 455031.384p 0.499711mV 455055.683p 0.476418mV 456035.002p 0.494899mV 456041.696p 0.475293mV 457005.969p 0.538178mV 458004.953p 0.575048mV 458015.406p 0.596021mV 458019.239p 0.596021mV 459000.836p 0.516831mV 459029.108p 0.493587mV 460028.662p 0.581731mV 461042.651p 0.61476mV 461044.751p 0.61476mV 461070.008p 0.773808mV 462023.178p 0.534087mV 462049.195p 0.46947mV 463020.723p 0.524988mV 463037.138p 0.46821mV 463045.04p 0.422191mV 463063.686p 0.338615mV 464002.321p 0.531021mV 464011.734p 0.525614mV 464022.361p 0.507098mV 464046.228p 0.465812mV 464051.925p 0.445126mV 465002.075p 0.548526mV 465030.805p 0.496989mV 465033.278p 0.496989mV 466014.925p 0.520037mV 466052.638p 0.362278mV 467031.089p 0.521745mV 467033.102p 0.521745mV 467045.12p 0.487892mV 467050.602p 0.467676mV 467052.871p 0.467676mV 468070.847p 0.3247mV 469004.411p 0.52613mV 469004.577p 0.52613mV 469012.476p 0.533969mV 469030.828p 0.598931mV 469035.493p 0.612252mV 469056.353p 0.681888mV 469064.114p 0.716353mV 469068.191p 0.757886mV 470006.921p 0.561582mV 470019.075p 0.57945mV 470050.628p 0.593722mV 470058.616p 0.594808mV 470065.989p 0.578926mV 470076.256p 0.551421mV 470080.988p 0.534683mV 470086.09p 0.524255mV 470122.536p 0.392474mV 470124.733p 0.392474mV 471002.065p 0.517383mV 471015.381p 0.512499mV 471028.63p 0.506026mV 471044.507p 0.478521mV 471068.241p 0.352335mV 472001.142p 0.566321mV 472030.278p 0.64048mV 472042.872p 0.6762mV 473057.4p 0.668107mV 474045.944p 0.421207mV 475001.03p 0.576215mV 475010.921p 0.583747mV 475059.06p 0.650763mV 475065.238p 0.678059mV 475073.443p 0.702119mV 475078.639p 0.733231mV 476013.441p 0.561223mV 476087.287p 0.633323mV 476111.048p 0.681259mV 476119.934p 0.701626mV 477006.896p 0.558377mV 477024.277p 0.571689mV 477029.148p 0.584702mV 477036.547p 0.617524mV 477074.559p 0.763105mV 478086.604p 0.479289mV 478110.802p 0.333219mV 479065.927p 0.425693mV 480023.211p 0.527611mV 480037.35p 0.505213mV 481013.814p 0.59949mV 481022.993p 0.605273mV 481031.24p 0.599749mV 481047.827p 0.571878mV 481059.797p 0.531282mV 481075.963p 0.436471mV 481078.707p 0.436471mV 481079.779p 0.436471mV 482017.673p 0.517278mV 482025.564p 0.534792mV 482040.384p 0.569441mV 482045.547p 0.593531mV 482050.829p 0.611442mV 482067.017p 0.692492mV 482079.55p 0.751947mV 483039.951p 0.614048mV 484026.743p 0.600069mV 484041.077p 0.618279mV 484044.014p 0.618279mV 484046.196p 0.620879mV 484074.475p 0.634628mV 484125.6p 0.710635mV 484149.483p 0.732142mV 484154.549p 0.743305mV 484155.871p 0.749409mV 484167.907p 0.759092mV 484169.928p 0.759092mV 484171.813p 0.762724mV 485007.192p 0.578111mV 485020.541p 0.577913mV 485022.242p 0.577913mV 485028.379p 0.578133mV 485045.097p 0.555398mV 485046.516p 0.555398mV 485067.34p 0.571584mV 485088.158p 0.577098mV 485124.083p 0.581998mV 486008.061p 0.515624mV 487010.895p 0.572239mV 487023.301p 0.603497mV 487043.05p 0.682126mV 487056.22p 0.748024mV 488049.018p 0.516002mV 488052.362p 0.498091mV 488054.926p 0.498091mV 488059.959p 0.486264mV 489003.807p 0.553124mV 489016.127p 0.548878mV 489016.463p 0.548878mV 489079.06p 0.581884mV 489082.183p 0.576624mV 489113.707p 0.566796mV 489119.329p 0.568545mV 489126.979p 0.591272mV 489197.072p 0.685843mV 489207.062p 0.722681mV 489217.165p 0.763326mV 490002.735p 0.601373mV 490068.417p 0.517451mV 490081.323p 0.516183mV 490092.883p 0.545649mV 490105.751p 0.63643mV 490111.327p 0.66708mV 491027.731p 0.506582mV 491029.34p 0.506582mV 492019.539p 0.534048mV 492023.584p 0.515427mV 492027.716p 0.490404mV 493008.572p 0.551698mV 493016.195p 0.571685mV 493057.763p 0.687032mV 493083.132p 0.762759mV 494027.438p 0.584172mV 494031.154p 0.578239mV 494054.201p 0.581607mV 494068.681p 0.642703mV 494071.417p 0.676322mV 494079.731p 0.716793mV 494080.136p 0.764297mV 495046.936p 0.473289mV 495052.421p 0.46361mV 495055.066p 0.459731mV 495055.068p 0.459731mV 495081.816p 0.475855mV 495132.692p 0.430385mV 496003.336p 0.597347mV 496028.915p 0.573414mV 496032.608p 0.56813mV 497027.543p 0.511855mV 497037.858p 0.493576mV 497038.17p 0.493576mV 497067.978p 0.442987mV 497080.893p 0.432406mV 497096.824p 0.408936mV 497105.15p 0.38711mV 497112.94p 0.384132mV 497114.477p 0.384132mV 497142.221p 0.400464mV 497182.187p 0.469009mV 497240.827p 0.586949mV 497247.006p 0.599989mV 497278.332p 0.680046mV 497286.038p 0.720108mV 497292.633p 0.732149mV 498001.209p 0.504854mV 498033.027p 0.457723mV 498052.736p 0.433265mV 498056.252p 0.44103mV 498067.681p 0.460661mV 498080.235p 0.476246mV 498087.394p 0.480479mV 498101.854p 0.452739mV 498115.417p 0.40125mV 499027.842p 0.527018mV 500011.611p 0.583165mV 500014.472p 0.583165mV 500024.855p 0.601763mV 500034.15p 0.634056mV 500044.546p 0.668011mV 500045.214p 0.695277mV 501002.754p 0.602955mV 502058.2p 0.577053mV 502064.395p 0.571753mV 502073.082p 0.58053mV 502081.295p 0.615126mV 502083.632p 0.615126mV 502089.924p 0.629653mV 502129.984p 0.703972mV 502136.635p 0.702494mV 502162.374p 0.744085mV 502168.373p 0.746973mV 502168.411p 0.746973mV 502177.128p 0.774962mV 503008.902p 0.548895mV 503028.892p 0.497469mV 503042.475p 0.41891mV 504012.808p 0.576383mV 504013.516p 0.576383mV 504035.962p 0.583227mV 504036.709p 0.583227mV 504048.758p 0.580886mV 504105.433p 0.4108mV 505002.734p 0.553967mV 505028.636p 0.489133mV 505037.195p 0.418131mV 506021.657p 0.561062mV 506046.635p 0.494607mV 506060.075p 0.452974mV 506064.093p 0.452974mV 506081.402p 0.402363mV 507001.97p 0.582716mV 507015.892p 0.603669mV 507029.796p 0.612608mV 507046.371p 0.61009mV 507074.793p 0.51142mV 507087.535p 0.404147mV 507088.316p 0.404147mV 507091.188p 0.363144mV 510007.538p 0.504264mV 510010.422p 0.5105mV 510015.686p 0.510152mV 510023.821p 0.503257mV 510050.851p 0.524869mV 510068.97p 0.560291mV 510097.133p 0.588026mV 510113.948p 0.58261mV 510128.346p 0.535184mV 510144.033p 0.53196mV 510165.45p 0.562016mV 510166.543p 0.562016mV 510183.981p 0.582413mV 510187.718p 0.581082mV 510221.298p 0.525824mV 510231.072p 0.493321mV 510269.135p 0.330554mV 511014.702p 0.50526mV 511020.199p 0.510805mV 511025.393p 0.522596mV 511061.065p 0.601521mV 511087.942p 0.73958mV 512017.083p 0.559122mV 512043.258p 0.527522mV 512096.913p 0.368116mV 512105.52p 0.370619mV 512136.816p 0.38864mV 512142.104p 0.390952mV 512179.355p 0.455777mV 512258.181p 0.467925mV 512286.713p 0.534907mV 512295.591p 0.592549mV 512314.762p 0.689584mV 512321.444p 0.763596mV 513026.826p 0.596079mV 513033.618p 0.603911mV 513042.283p 0.614197mV 513042.454p 0.614197mV 513053.33p 0.651095mV 513063.311p 0.702607mV 513069.158p 0.732604mV 514031.345p 0.464463mV 515016.163p 0.539236mV 515016.567p 0.539236mV 515018.04p 0.539236mV 515047.98p 0.656743mV 515048.963p 0.656743mV 515054.395p 0.676566mV 516001.871p 0.519167mV 516072.127p 0.388392mV 516078.571p 0.380682mV 516099.391p 0.364275mV 516113.017p 0.346564mV 516124.253p 0.343095mV 516167.063p 0.387461mV 516186.762p 0.337777mV 517008.451p 0.554618mV 517026.333p 0.568183mV 517036.325p 0.600349mV 517044.099p 0.619871mV 518002.408p 0.556702mV 518005.144p 0.556767mV 518047.53p 0.701677mV 519013.538p 0.564895mV 519018.822p 0.565498mV 519047.383p 0.513933mV 519055.159p 0.496329mV 519093.348p 0.476811mV 520015.672p 0.509479mV 520065.838p 0.481125mV 520080.758p 0.454935mV 520099.305p 0.41752mV 521010.767p 0.535089mV 521016.427p 0.535028mV 521022.311p 0.528573mV 521026.63p 0.528324mV 521028.487p 0.528324mV 522017.014p 0.562682mV 523011.862p 0.543924mV 523024.84p 0.513062mV 523055.814p 0.48903mV 523058.945p 0.48903mV 523060.498p 0.480649mV 523062.543p 0.480649mV 524009.949p 0.580307mV 524036.193p 0.712297mV 525006.623p 0.564567mV 525019.007p 0.556431mV 525055.527p 0.718642mV 525064.739p 0.752054mV 526032.382p 0.572003mV 526032.64p 0.572003mV 526042.312p 0.57958mV 526046.467p 0.580431mV 526058.805p 0.576398mV 526060.207p 0.571485mV 526064.22p 0.571485mV 526064.909p 0.571485mV 526070.764p 0.54323mV 526101.239p 0.50794mV 527007.992p 0.521303mV 527034.273p 0.617738mV 527045.912p 0.727951mV 527051.24p 0.761967mV 528016.735p 0.575547mV 528018.835p 0.575547mV 528021.284p 0.581637mV 528048.357p 0.595874mV 528061.14p 0.599442mV 528112.416p 0.630548mV 528117.084p 0.624416mV 528121.989p 0.612509mV 528149.748p 0.514215mV 529004.038p 0.557866mV 529010.006p 0.56298mV 529023.992p 0.580919mV 529028.514p 0.580638mV 529039.413p 0.599555mV 529041.07p 0.618789mV 529045.038p 0.644628mV 530015.101p 0.604931mV 530029.04p 0.613768mV 531008.994p 0.543183mV 531046.877p 0.524865mV 531100.011p 0.651449mV 531107.211p 0.676933mV 532011.052p 0.513162mV 532023.918p 0.506278mV 532068.345p 0.36955mV 532164.353p 0.519454mV 532195.627p 0.663429mV 533001.827p 0.556471mV 533025.467p 0.535656mV 533025.679p 0.535656mV 533054.965p 0.55733mV 533055.227p 0.557684mV 533093.354p 0.420293mV 534003.218p 0.50714mV 534021.269p 0.527929mV 534049.279p 0.607248mV 535034.624p 0.527896mV 535090.831p 0.520025mV 535091.87p 0.520025mV 535121.431p 0.592073mV 535136.674p 0.664229mV 536004.968p 0.53846mV 536012.418p 0.546327mV 536025.48p 0.541997mV 536039.368p 0.536809mV 536087.619p 0.501377mV 536093.781p 0.493307mV 536122.496p 0.417479mV 536127.734p 0.387184mV 537019.67p 0.560541mV 537052.077p 0.509154mV 537057.569p 0.508555mV 537074.282p 0.505232mV 538015.456p 0.575727mV 538054.4p 0.513841mV 539013.214p 0.555036mV 539015.59p 0.554197mV 539017.972p 0.554197mV 539062.661p 0.434331mV 539080.759p 0.340146mV 540000.986p 0.500477mV 540102.678p 0.526804mV 540118.642p 0.518736mV 540124.063p 0.507316mV 540135.648p 0.471633mV 541013.061p 0.501814mV 541063.149p 0.442001mV 541093.136p 0.388034mV 541105.404p 0.339286mV 542011.335p 0.585471mV 542039.409p 0.57688mV 542053.334p 0.582041mV 542058.694p 0.584061mV 542066.814p 0.59502mV 542076.131p 0.619605mV 542077.775p 0.619605mV 543011.322p 0.518504mV 543014.549p 0.518504mV 543057.083p 0.553024mV 543060.354p 0.569546mV 543083.915p 0.624136mV 543107.915p 0.698239mV 543110.415p 0.706434mV 543123.505p 0.706974mV 543137.412p 0.680938mV 544017.139p 0.502479mV 544044.505p 0.515236mV 544047.695p 0.513101mV 544048.201p 0.513101mV 544065.41p 0.48951mV 544069.531p 0.48951mV 544092.657p 0.461269mV 544127.77p 0.37658mV 545003.791p 0.546743mV 545120.917p 0.3489mV 545124.805p 0.3489mV 546000.287p 0.552776mV 546017.847p 0.574865mV 546029.099p 0.621438mV 546030.392p 0.641938mV 546048.498p 0.719244mV 546052.426p 0.742419mV 546054.842p 0.742419mV 547011.479p 0.516647mV 547024.994p 0.522724mV 547047.212p 0.60794mV 547048.856p 0.60794mV 547051.175p 0.639067mV 548002.753p 0.582351mV 548019.561p 0.586611mV 548066.909p 0.516143mV 548074.326p 0.533803mV 548084.643p 0.549698mV 548144.785p 0.73467mV 549029.264p 0.573965mV 549040.51p 0.60533mV 549062.36p 0.579863mV 549102.883p 0.474343mV 550000.474p 0.517255mV 550001.598p 0.517255mV 550034.599p 0.535232mV 550037.753p 0.546992mV 550060.493p 0.68838mV 551009.029p 0.57302mV 551020.889p 0.572716mV 551025.416p 0.585437mV 551029.143p 0.585437mV 551068.179p 0.748383mV 552002.852p 0.549266mV 552019.93p 0.542683mV 552044.366p 0.59872mV 552067.307p 0.742951mV 553006.144p 0.521921mV 553017.914p 0.52972mV 553059.831p 0.518939mV 553079.501p 0.491338mV 553083.154p 0.471214mV 554001.256p 0.583855mV 554013.246p 0.576668mV 554019.909p 0.563943mV 554020.192p 0.545088mV 554043.75p 0.406168mV 554046.952p 0.367267mV 555017.438p 0.607581mV 555030.333p 0.661762mV 555046.642p 0.727596mV 556002.813p 0.533329mV 556004.697p 0.533329mV 556018.968p 0.541297mV 556025.202p 0.535731mV 556050.422p 0.593313mV 556052.349p 0.593313mV 556067.351p 0.677299mV 556068.922p 0.677299mV 557016.879p 0.531361mV 557037.074p 0.552695mV 557041.556p 0.557974mV 557045.36p 0.556969mV 557049.308p 0.556969mV 557058.284p 0.574007mV 557072.371p 0.647681mV 557075.074p 0.685466mV 557084.778p 0.730131mV 558001.944p 0.50844mV 558010.375p 0.514679mV 558022.61p 0.532502mV 558071.056p 0.663706mV 558088.921p 0.741572mV 559002.562p 0.569351mV 559054.705p 0.573324mV 559062.545p 0.570445mV 559090.754p 0.514388mV 560000.137p 0.508424mV 560004.758p 0.508424mV 560013.919p 0.513674mV 560018.15p 0.525347mV 560062.346p 0.673881mV 560077.332p 0.747587mV 561004.258p 0.547497mV 561006.538p 0.547488mV 561022.376p 0.560008mV 561023.587p 0.560008mV 561038.719p 0.617009mV 561055.236p 0.684931mV 561065.12p 0.710403mV 562065.283p 0.612246mV 562072.633p 0.62914mV 562072.924p 0.62914mV 562075.58p 0.652714mV 562090.068p 0.726917mV 563027.438p 0.545249mV 563032.159p 0.550091mV 563037.593p 0.561205mV 563059.872p 0.543155mV 563085.878p 0.465374mV 563089.462p 0.465374mV 564002.398p 0.568571mV 564035.478p 0.570899mV 564059.347p 0.646249mV 564073.307p 0.700965mV 565049.66p 0.424863mV 566020.382p 0.540073mV 566032.826p 0.59627mV 566053.692p 0.686055mV 566060.504p 0.747179mV 566063.626p 0.747179mV 567004.072p 0.597688mV 567015.569p 0.593121mV 567082.091p 0.488953mV 567138.364p 0.501207mV 567151.934p 0.502215mV 567153.866p 0.502215mV 567169.264p 0.519422mV 567179.225p 0.514992mV 567179.734p 0.514992mV 567181.319p 0.503045mV 568022.217p 0.578177mV 568034.347p 0.598664mV 568050.203p 0.668433mV 568053.336p 0.668433mV 569002.489p 0.562216mV 569005.348p 0.561885mV 569011.528p 0.567934mV 569018.279p 0.580358mV 569038.517p 0.644437mV 569057.073p 0.703373mV 569058.013p 0.703373mV 569061.819p 0.71383mV 570025.329p 0.530284mV 570037.32p 0.487191mV 570043.107p 0.468491mV 571004.34p 0.549596mV 571026.868p 0.51883mV 571027.352p 0.51883mV 571035.287p 0.496831mV 571064.57p 0.388909mV 572027.12p 0.539952mV 572045.018p 0.539671mV 572067.792p 0.47495mV 573001.162p 0.503818mV 573001.31p 0.503818mV 573011.535p 0.511862mV 573015.459p 0.524897mV 573043.83p 0.568923mV 574013.641p 0.549158mV 574057.833p 0.500153mV 574073.496p 0.520523mV 574122.894p 0.629166mV 574138.782p 0.695192mV 575006.36p 0.506061mV 575008.376p 0.506061mV 575009.016p 0.506061mV 575033.441p 0.462324mV 575051.626p 0.328522mV 576012.786p 0.553002mV 576017.548p 0.564888mV 576037.322p 0.55016mV 576038.93p 0.55016mV 576120.022p 0.480161mV 576140.292p 0.497573mV 576146.319p 0.513482mV 576174.019p 0.545694mV 576179.116p 0.548178mV 576192.9p 0.555489mV 576204.317p 0.566604mV 576212.299p 0.590561mV 576216.138p 0.60594mV 576217.594p 0.60594mV 576217.741p 0.60594mV 576233.333p 0.65394mV 576238.048p 0.683412mV 576242.22p 0.707264mV 577005.006p 0.554442mV 577008.364p 0.554442mV 577031.75p 0.61513mV 577044.567p 0.637194mV 577090.971p 0.698298mV 577099.671p 0.708273mV 577116.69p 0.733108mV 577121.459p 0.729627mV 577124.87p 0.729627mV 577125.432p 0.73349mV 577131.157p 0.732278mV 577133.511p 0.732278mV 577142.417p 0.751889mV 577142.759p 0.751889mV 577150.896p 0.763901mV 577152.126p 0.763901mV 577152.602p 0.763901mV 578007.601p 0.599817mV 578028.462p 0.591834mV 578036.34p 0.589476mV 578045.848p 0.613289mV 578058.526p 0.638353mV 578066.415p 0.690419mV 579002.532p 0.538114mV 579010.197p 0.533298mV 579023.093p 0.515557mV 579027.217p 0.515903mV 579062.958p 0.576929mV 579067.483p 0.601689mV 579074.74p 0.632916mV 580022.314p 0.517295mV 580059.402p 0.576299mV 580064.657p 0.605888mV 580076.384p 0.65858mV 580088.754p 0.665127mV 580094.775p 0.660071mV 580120.166p 0.624915mV 580143.735p 0.637788mV 580157.426p 0.680912mV 580161.603p 0.696675mV 581010.921p 0.551992mV 581020.816p 0.569402mV 581027.151p 0.568748mV 581053.221p 0.611866mV 581064.087p 0.632337mV 581080.382p 0.692044mV 581093.05p 0.720152mV 581094.755p 0.720152mV 581104.07p 0.7522mV 581108.816p 0.760639mV 582001.006p 0.594946mV 582024.249p 0.638731mV 582051.483p 0.694889mV 582074.331p 0.765908mV 583035.373p 0.561368mV 583048.061p 0.603845mV 583057.99p 0.647097mV 584012.415p 0.595754mV 584061.966p 0.615004mV 585003.166p 0.538364mV 585018.179p 0.520928mV 585023.62p 0.502336mV 585042.041p 0.437693mV 585051.266p 0.414765mV 585054.704p 0.414765mV 586027.995p 0.479782mV 586047.182p 0.356311mV 586049.357p 0.356311mV 587026.401p 0.530379mV 587077.247p 0.493096mV 587095.537p 0.458423mV 587104.227p 0.448532mV 587155.694p 0.39044mV 588027.966p 0.495422mV 588064.793p 0.354078mV 589013.521p 0.518078mV 589049.918p 0.449948mV 590011.033p 0.525406mV 590035.541p 0.445112mV 591040.139p 0.550286mV 591045.321p 0.536834mV 591051.019p 0.529686mV 591090.498p 0.531669mV 591095.027p 0.529825mV 591097.113p 0.529825mV 591151.126p 0.458979mV 591152.538p 0.458979mV 592010.213p 0.550465mV 592013.232p 0.550465mV 593012.632p 0.589612mV 593019.767p 0.589973mV 593036.859p 0.631923mV 593061.725p 0.754913mV 594015.644p 0.594016mV 594019.127p 0.594016mV 594029.632p 0.603524mV 594046.231p 0.664431mV 594052.768p 0.674651mV 595072.211p 0.4646mV 595101.653p 0.404198mV 596011.319p 0.602694mV 596045.272p 0.646397mV 596082.217p 0.747427mV 596082.516p 0.747427mV 596086.116p 0.768956mV 597008.701p 0.498122mV 597051.422p 0.547312mV 597060.437p 0.547904mV 597089.009p 0.571587mV 597095.257p 0.560407mV 597117.45p 0.539094mV 597146.339p 0.454119mV 598009.045p 0.512714mV 598009.868p 0.512714mV 598075.84p 0.622823mV 598086.035p 0.690151mV 599001.376p 0.540592mV 599007.799p 0.540096mV 599034.402p 0.492271mV 599072.351p 0.532588mV 599075.272p 0.553193mV 599097.46p 0.597806mV 599104.685p 0.612535mV 599114.777p 0.661867mV 599124.235p 0.738448mV 600057.568p 0.431032mV 600085.635p 0.381847mV 601016.561p 0.558956mV 601087.51p 0.611726mV 603004.211p 0.577245mV 603024.466p 0.577106mV 603030.497p 0.584217mV 603046.53p 0.618436mV 603056.785p 0.653401mV 603072.524p 0.738435mV 604005.587p 0.501246mV 604013.817p 0.507414mV 604036.568p 0.451956mV 605001.14p 0.585811mV 605020.928p 0.548559mV 605031.005p 0.530761mV 605055.708p 0.544371mV 605058.027p 0.544371mV 605069.434p 0.575433mV 605113.851p 0.603261mV 605117.101p 0.593586mV 605121.098p 0.577954mV 605136.408p 0.494484mV 605136.439p 0.494484mV 606007.658p 0.561316mV 606014.502p 0.554824mV 606029.254p 0.535652mV 606031.68p 0.52928mV 606038.481p 0.529119mV 606071.161p 0.627755mV 606073.944p 0.627755mV 606076.882p 0.640994mV 606097.926p 0.67446mV 606103.265p 0.672055mV 606111.876p 0.663326mV 606161.414p 0.765686mV 606164.61p 0.765686mV 607022.553p 0.520769mV 607030.485p 0.462302mV 608000.461p 0.519677mV 608019.952p 0.539712mV 608026.823p 0.558634mV 608034.616p 0.564886mV 608046.594p 0.621975mV 608114.461p 0.708715mV 608119.993p 0.710096mV 608128.822p 0.734523mV 608133.114p 0.745192mV 608138.02p 0.75082mV 609033.192p 0.512728mV 609037.392p 0.500096mV 609041.494p 0.493528mV 609050.778p 0.460526mV 610006.122p 0.600809mV 610013.507p 0.595815mV 610119.924p 0.409643mV 611011.485p 0.552076mV 611015.194p 0.539849mV 612033.878p 0.580289mV 612044.85p 0.616369mV 612048.657p 0.631642mV 612072.37p 0.760732mV 613009.23p 0.554333mV 613033.009p 0.62177mV 613064.974p 0.714134mV 613071.442p 0.755587mV 614023.318p 0.544345mV 614055.782p 0.677131mV 616002.38p 0.537575mV 616069.884p 0.488484mV 616085.416p 0.534301mV 616118.32p 0.688698mV 616137.982p 0.745291mV 616149.969p 0.75525mV 616151.502p 0.752843mV 617002.497p 0.578991mV 617005.221p 0.578298mV 617023.056p 0.602536mV 617068.463p 0.615089mV 617094.871p 0.716324mV 618013.055p 0.517855mV 618021.383p 0.521152mV 618042.57p 0.512798mV 618061.148p 0.488551mV 618063.003p 0.488551mV 618122.694p 0.325715mV 619012.143p 0.515071mV 619028.699p 0.568304mV 619059.459p 0.747295mV 620020.658p 0.591608mV 620021.891p 0.591608mV 620040.067p 0.644665mV 620067.712p 0.697754mV 621030.377p 0.562047mV 621037.803p 0.562744mV 621081.46p 0.449353mV 621091.599p 0.366448mV 622017.013p 0.604852mV 622017.932p 0.604852mV 622028.275p 0.599171mV 622034.971p 0.593662mV 622083.697p 0.399917mV 623061.181p 0.57593mV 623066.127p 0.585296mV 623074.18p 0.601126mV 623088.482p 0.61254mV 623089.155p 0.61254mV 623120.893p 0.595537mV 623167.253p 0.4673mV 624010.426p 0.548492mV 624012.648p 0.548492mV 624042.287p 0.560725mV 624070.542p 0.523143mV 625036.664p 0.527546mV 625042.406p 0.496599mV 625044.344p 0.496599mV 625054.174p 0.440395mV 625069.341p 0.342321mV 626008.775p 0.555221mV 626042.174p 0.511603mV 626048.828p 0.485488mV 626049.419p 0.485488mV 627004.712p 0.575667mV 627032.753p 0.565433mV 627034.361p 0.565433mV 627105.137p 0.430875mV 627123.498p 0.415177mV 627124.651p 0.415177mV 627126.924p 0.420799mV 627134.673p 0.419329mV 627156.883p 0.40557mV 627165.56p 0.38511mV 627196.364p 0.373819mV 628016.033p 0.516821mV 628026.419p 0.536215mV 628041.398p 0.598996mV 628049.919p 0.611706mV 628057.275p 0.644428mV 628066.895p 0.691697mV 629007.567p 0.580889mV 629014.318p 0.587644mV 629048.859p 0.680551mV 629054.075p 0.703018mV 630019.118p 0.53777mV 630024.266p 0.531928mV 630039.112p 0.475948mV 630040.727p 0.444223mV 630043.534p 0.444223mV 631022.387p 0.587167mV 631031.865p 0.583868mV 631048.997p 0.53334mV 632000.4p 0.581054mV 632002.321p 0.581054mV 632014.77p 0.573092mV 632022.301p 0.565849mV 632030.506p 0.546538mV 632038.683p 0.546403mV 632051.894p 0.571111mV 632079.28p 0.635779mV 632105.525p 0.595964mV 632126.116p 0.578284mV 632129.564p 0.578284mV 632130.091p 0.590044mV 632133.773p 0.590044mV 632140.186p 0.620473mV 632140.262p 0.620473mV 632154.977p 0.652331mV 632158.478p 0.672176mV 632161.389p 0.698932mV 632172.989p 0.77364mV 633014.437p 0.531116mV 633032.04p 0.590014mV 633032.872p 0.590014mV 633037.602p 0.601725mV 633050.428p 0.663896mV 634021.717p 0.49647mV 634053.685p 0.389588mV 634067.449p 0.390642mV 635018.122p 0.531516mV 635020.297p 0.538296mV 635024.357p 0.538296mV 635074.829p 0.736921mV 636023.845p 0.573666mV 636036.718p 0.63307mV 637003.847p 0.585601mV 637019.409p 0.576945mV 637041.074p 0.659147mV 637056.382p 0.696597mV 637064.401p 0.706481mV 637120.008p 0.757016mV 638004.228p 0.522058mV 638004.547p 0.522058mV 638022.307p 0.53343mV 638044.888p 0.606016mV 638053.25p 0.63688mV 638057.253p 0.66235mV 638060.078p 0.694641mV 640000.226p 0.555027mV 640002.517p 0.555027mV 640037.8p 0.482475mV 640048.211p 0.460636mV 640067.821p 0.334984mV 641007.031p 0.547379mV 641042.994p 0.451569mV 641080.593p 0.465656mV 641085.575p 0.472313mV 641121.039p 0.41574mV 641128.366p 0.417416mV 641138.841p 0.399508mV 642114.997p 0.650461mV 642132.975p 0.700147mV 642132.977p 0.700147mV 642133.209p 0.700147mV 642140.275p 0.742062mV 642146.393p 0.773865mV 643008.311p 0.516963mV 643010.247p 0.511022mV 643015.976p 0.498575mV 643018.78p 0.498575mV 643026.07p 0.453978mV 643029.292p 0.453978mV 644012.001p 0.562671mV 644031.742p 0.566356mV 644048.648p 0.589227mV 644062.522p 0.607395mV 644072.233p 0.606362mV 644083.888p 0.59422mV 644105.182p 0.591176mV 644113.147p 0.590219mV 644124.424p 0.57019mV 644130.962p 0.56356mV 644131.547p 0.56356mV 644133.918p 0.56356mV 644141.293p 0.557315mV 644167.249p 0.602755mV 644184.84p 0.637378mV 644202.16p 0.648541mV 644218.994p 0.663343mV 644228.678p 0.657893mV 644241.984p 0.664295mV 644253.383p 0.665918mV 644285.788p 0.71098mV 644289.64p 0.71098mV 645002.664p 0.570103mV 645014.555p 0.577052mV 645028.281p 0.610694mV 645054.553p 0.703207mV 645064.451p 0.756278mV 646006.146p 0.531863mV 646007.706p 0.531863mV 646015.224p 0.525756mV 646057.938p 0.649899mV 647027.282p 0.563221mV 647035.153p 0.567441mV 647038.88p 0.567441mV 647071.227p 0.511324mV 647080.867p 0.515032mV 647106.291p 0.466395mV 648047.718p 0.686755mV 649008.498p 0.575952mV 649019.408p 0.583806mV 649053.197p 0.518072mV 649058.956p 0.519304mV 649059.216p 0.519304mV 649062.066p 0.514035mV 649107.779p 0.551209mV 649110.168p 0.569209mV 649152.422p 0.69556mV 649159.605p 0.710634mV 649162.814p 0.720385mV 649188.787p 0.767231mV 650015.355p 0.578546mV 650026.982p 0.587742mV 650049.925p 0.621682mV 650054.096p 0.618513mV 650066.23p 0.586459mV 650070.003p 0.572251mV 650076.331p 0.551976mV 650083.533p 0.52554mV 650089.561p 0.492814mV 651001.942p 0.520635mV 651007.737p 0.521445mV 651030.961p 0.4915mV 652005.195p 0.592315mV 652020.293p 0.596269mV 652029.41p 0.585617mV 652069.231p 0.377231mV 653017.101p 0.546653mV 653027.191p 0.554631mV 653030.36p 0.561784mV 653045.117p 0.621446mV 653049.738p 0.621446mV 653050.647p 0.641752mV 653067.281p 0.743568mV 654001.233p 0.542615mV 654014.484p 0.534397mV 654016.087p 0.520759mV 654052.948p 0.379991mV 655001.48p 0.521493mV 655003.484p 0.521493mV 655012.097p 0.526827mV 655012.445p 0.526827mV 655036.519p 0.534017mV 656018.04p 0.493213mV 656038.533p 0.423806mV 657026.785p 0.549002mV 657049.081p 0.609791mV 657055.612p 0.616364mV 657091.331p 0.720564mV 658051.388p 0.592518mV 658068.642p 0.627506mV 658091.684p 0.737699mV 658094.555p 0.737699mV 659002.097p 0.575181mV 659015.926p 0.558499mV 659043.136p 0.455825mV 659048.78p 0.443218mV 659113.065p 0.506324mV 659118.082p 0.534136mV 659129.539p 0.608009mV 659140.407p 0.755028mV 660018.304p 0.520014mV 660026.236p 0.538914mV 660038.308p 0.557259mV 660051.964p 0.594284mV 660089.79p 0.544542mV 661063.611p 0.612216mV 661066.408p 0.602636mV 661071.367p 0.587158mV 661072.494p 0.587158mV 661076.247p 0.565718mV 662020.856p 0.503145mV 662025.811p 0.502053mV 662032.072p 0.494371mV 662068.605p 0.519759mV 662099.043p 0.590077mV 662106.872p 0.639057mV 663007.756p 0.499529mV 664036.01p 0.73228mV 665015.643p 0.508851mV 665049.331p 0.449964mV 665049.757p 0.449964mV 665094.367p 0.575143mV 665095.485p 0.592709mV 665103.855p 0.604134mV 665135.222p 0.630491mV 665158.229p 0.691051mV 665181.001p 0.710029mV 665181.378p 0.710029mV 665185.93p 0.700633mV 665186.569p 0.700633mV 665187.223p 0.700633mV 665210.258p 0.623672mV 665224.084p 0.584004mV 666003.544p 0.579264mV 666011.957p 0.586087mV 666014.799p 0.586087mV 666049.025p 0.575399mV 666085.287p 0.712424mV 666096.938p 0.768411mV 667000.224p 0.541691mV 667011.685p 0.533394mV 667017.899p 0.519709mV 667036.829p 0.399895mV 667036.92p 0.399895mV 667044.781p 0.365524mV 668015.25p 0.548514mV 668019.228p 0.548514mV 668031.228p 0.523952mV 668041.31p 0.530194mV 668042.842p 0.530194mV 668055.276p 0.57317mV 668061.109p 0.591692mV 668062.662p 0.591692mV 668064.177p 0.591692mV 668065.003p 0.60406mV 668067.163p 0.60406mV 668077.701p 0.610777mV 668109.673p 0.665837mV 668118.192p 0.680291mV 668121.435p 0.691795mV 668122.392p 0.691795mV 668122.44p 0.691795mV 668130.049p 0.723588mV 668130.105p 0.723588mV 668138.567p 0.731592mV 668148.317p 0.732296mV 668150.703p 0.73747mV 668154.736p 0.73747mV 668155.992p 0.749985mV 668177.644p 0.775261mV 669007.147p 0.567842mV 669033.02p 0.565161mV 669052.712p 0.481719mV 670010.616p 0.533163mV 670016.639p 0.545415mV 670034.121p 0.607086mV 670038.469p 0.632131mV 670046.064p 0.689751mV 670064.778p 0.734927mV 670065.729p 0.739607mV 670082.88p 0.735907mV 671001.592p 0.519449mV 671052.034p 0.522486mV 671055.898p 0.508536mV 671058.913p 0.508536mV 671064.312p 0.500712mV 671119.862p 0.482097mV 671143.157p 0.59489mV 671150.15p 0.63382mV 671155.066p 0.650667mV 671160.753p 0.661761mV 671190.518p 0.763167mV 672007.94p 0.566798mV 672024.186p 0.552111mV 672026.065p 0.538947mV 672040.223p 0.461355mV 672054.803p 0.376613mV 673000.952p 0.595395mV 673009.355p 0.595245mV 673033.718p 0.630801mV 673034.375p 0.630801mV 673050.442p 0.667645mV 673053.074p 0.667645mV 673053.176p 0.667645mV 673071.192p 0.740865mV 674000.341p 0.501542mV 674045.349p 0.587396mV 674068.506p 0.699104mV 674069.742p 0.699104mV 674072.937p 0.731625mV 675011.863p 0.598553mV 675012.809p 0.598553mV 675046.494p 0.558936mV 675054.493p 0.55601mV 675055.858p 0.546839mV 675083.935p 0.443069mV 676036.097p 0.633109mV 676073.36p 0.672868mV 676127.119p 0.598324mV 676153.906p 0.619886mV 676197.841p 0.771562mV 677023.402p 0.56269mV 677037.843p 0.617768mV 677044.028p 0.624068mV 677058.786p 0.633077mV 677069.247p 0.656225mV 677082.173p 0.704901mV 677087.605p 0.72267mV 678013.597p 0.539803mV 678025.89p 0.534863mV 678106.41p 0.356554mV 678119.417p 0.355253mV 678126.997p 0.349067mV 678149.761p 0.333893mV 679006.44p 0.595706mV 679009.621p 0.595706mV 679021.896p 0.598389mV 679029.042p 0.599806mV 679035.921p 0.597269mV 679042.228p 0.593294mV 679044.839p 0.593294mV 679067.163p 0.621999mV 680045.653p 0.510488mV 680048.223p 0.510488mV 680084.512p 0.461096mV 680109.515p 0.437264mV 680109.691p 0.437264mV 680144.24p 0.411641mV 680149.234p 0.424068mV 680176.84p 0.590677mV 680193.351p 0.694221mV 680198.861p 0.717332mV 681005.09p 0.517914mV 681007.423p 0.517914mV 681038.123p 0.42392mV 682019.767p 0.560191mV 682022.274p 0.554124mV 682028.9p 0.554422mV 682037.31p 0.5614mV 682087.475p 0.602401mV 682105.289p 0.625288mV 682122.792p 0.649647mV 682134.124p 0.65402mV 682140.766p 0.673526mV 682151.083p 0.720896mV 683039.251p 0.467536mV 683051.3p 0.384878mV 684008.426p 0.5821mV 684011.605p 0.576224mV 684024.847p 0.558745mV 684047.467p 0.525371mV 684077.212p 0.405701mV 685001.033p 0.575105mV 685019.771p 0.569363mV 685037.323p 0.584685mV 685050.283p 0.57611mV 685061.333p 0.560844mV 685064.835p 0.560844mV 685065.893p 0.56284mV 685070.624p 0.558603mV 685088.99p 0.508423mV 685090.98p 0.491589mV 685096.896p 0.480791mV 685110.182p 0.445854mV 685126.854p 0.424422mV 685231.43p 0.462779mV 685292.193p 0.414107mV 686017.614p 0.560568mV 686026.482p 0.579259mV 686029.933p 0.579259mV 686030.39p 0.585592mV 686071.069p 0.713403mV 687007.882p 0.56042mV 687045.406p 0.579958mV 687053.02p 0.600086mV 687060.733p 0.647336mV 687077.444p 0.700043mV 687090.0p 0.728717mV 687093.501p 0.753868mV 688017.485p 0.548518mV 688086.607p 0.752887mV 689025.214p 0.619877mV 689052.39p 0.747341mV 690014.978p 0.512412mV 690022.153p 0.542543mV 690026.907p 0.566777mV 690054.168p 0.607804mV 690103.715p 0.646405mV 690128.95p 0.587347mV 690166.603p 0.415682mV 691001.351p 0.584286mV 691053.418p 0.429005mV 692029.661p 0.470286mV 692052.658p 0.367674mV 693041.698p 0.69948mV 694008.706p 0.60035mV 694021.364p 0.628791mV 694024.57p 0.628791mV 694053.466p 0.768952mV 695016.817p 0.588032mV 695032.985p 0.605576mV 695061.05p 0.644391mV 695066.83p 0.649463mV 695075.052p 0.680238mV 695080.833p 0.706036mV 695086.641p 0.738897mV 696031.549p 0.54745mV 696050.925p 0.580988mV 696071.347p 0.666981mV 697025.477p 0.488192mV 697031.7p 0.480477mV 697035.548p 0.478662mV 697040.012p 0.470122mV 697074.814p 0.374991mV 698001.644p 0.566999mV 698016.125p 0.583093mV 698028.899p 0.61341mV 698032.424p 0.632139mV 698052.453p 0.661763mV 698058.078p 0.676993mV 699013.405p 0.535534mV 699033.789p 0.6266mV 699039.564p 0.665452mV 700000.296p 0.568295mV 700010.272p 0.573921mV 700029.843p 0.592772mV 700039.192p 0.637781mV 701016.697p 0.58436mV 701016.879p 0.58436mV 701046.594p 0.564163mV 701073.841p 0.583092mV 701089.904p 0.586727mV 701107.272p 0.590462mV 701120.101p 0.617856mV 701124.518p 0.617856mV 701141.607p 0.73129mV 701142.717p 0.73129mV 702014.803p 0.543848mV 702018.47p 0.555622mV 702028.127p 0.585429mV 702053.877p 0.552952mV 702055.752p 0.540772mV 702092.284p 0.362389mV 703070.631p 0.454562mV 704020.318p 0.501247mV 704036.552p 0.513795mV 704042.853p 0.529959mV 704051.883p 0.568001mV 704063.403p 0.580854mV 704070.2p 0.606959mV 704084.209p 0.634126mV 704085.01p 0.657745mV 704098.519p 0.700419mV 704098.534p 0.700419mV 704100.12p 0.719759mV 704103.272p 0.719759mV 705008.378p 0.533082mV 705014.949p 0.539473mV 705018.211p 0.539457mV 705032.117p 0.513762mV 705044.19p 0.493742mV 705066.784p 0.49787mV 705151.041p 0.514183mV 705151.745p 0.514183mV 705154.878p 0.514183mV 705182.74p 0.446003mV 705196.143p 0.44489mV 705206.679p 0.45953mV 705210.314p 0.456517mV 705246.032p 0.380183mV 705254.936p 0.346624mV 706018.089p 0.510012mV 706064.676p 0.504313mV 706070.888p 0.479987mV 706087.095p 0.475174mV 706095.57p 0.459216mV 706107.631p 0.466253mV 706123.182p 0.469529mV 706135.838p 0.436738mV 707050.481p 0.477536mV 707051.616p 0.477536mV 707086.71p 0.341742mV 708002.307p 0.591757mV 708042.954p 0.539092mV 708077.591p 0.492066mV 708078.156p 0.492066mV 708097.348p 0.540992mV 708105.987p 0.557955mV 708111.271p 0.575837mV 708116.75p 0.600071mV 708130.055p 0.649118mV 708140.291p 0.694705mV 708142.028p 0.694705mV 708158.287p 0.747254mV 709040.936p 0.668445mV 709053.044p 0.705752mV 710029.523p 0.535mV 710033.177p 0.539338mV 710079.955p 0.598237mV 710104.171p 0.564787mV 710131.055p 0.586106mV 710209.379p 0.332542mV 711029.703p 0.600531mV 711050.317p 0.53954mV 711077.354p 0.371315mV 712028.577p 0.469439mV 712070.875p 0.434483mV 712083.623p 0.473294mV 712095.937p 0.511513mV 712101.646p 0.519307mV 712126.163p 0.574304mV 712133.785p 0.58135mV 712198.492p 0.557943mV 712209.938p 0.549502mV 712215.32p 0.528592mV 712218.889p 0.528592mV 712223.76p 0.514896mV 712241.806p 0.445177mV 712252.208p 0.432523mV 713000.835p 0.594993mV 713031.987p 0.507875mV 713041.518p 0.441518mV 713051.269p 0.398369mV 713065.332p 0.336657mV 714000.151p 0.56092mV 714004.402p 0.56092mV 714010.922p 0.565623mV 714014.905p 0.565623mV 714057.437p 0.535042mV 714100.819p 0.335622mV 715008.878p 0.600583mV 715043.243p 0.627361mV 715049.592p 0.653912mV 715050.953p 0.674664mV 715056.609p 0.702335mV 716009.498p 0.550198mV 716032.049p 0.489265mV 716055.009p 0.363703mV 717040.851p 0.628637mV 717058.768p 0.687026mV 718007.605p 0.581644mV 718021.304p 0.572381mV 718031.123p 0.543948mV 718031.315p 0.543948mV 718051.939p 0.436385mV 718067.346p 0.378897mV 718078.76p 0.354635mV 719001.068p 0.580441mV 719003.138p 0.580441mV 719031.74p 0.644596mV 719038.39p 0.647229mV 719047.68p 0.63548mV 719082.576p 0.627631mV 719121.904p 0.746988mV 720015.063p 0.531297mV 720072.7p 0.664188mV 720089.13p 0.724847mV 721020.993p 0.595683mV 721038.422p 0.620296mV 721048.898p 0.669894mV 722029.345p 0.528908mV 723002.216p 0.583485mV 723003.996p 0.583485mV 723021.172p 0.613818mV 724002.409p 0.551731mV 724014.071p 0.559865mV 724016.468p 0.573407mV 724065.758p 0.731749mV 725003.93p 0.524218mV 725013.661p 0.51766mV 725021.183p 0.51041mV 725027.546p 0.49703mV 725047.41p 0.440031mV 725047.49p 0.440031mV 725067.711p 0.436091mV 726013.033p 0.568155mV 726016.563p 0.555439mV 726046.784p 0.408134mV 727012.072p 0.584726mV 727018.852p 0.584592mV 727032.06p 0.572865mV 727073.959p 0.684448mV 727081.743p 0.760545mV 728019.951p 0.499168mV 728020.465p 0.504371mV 728032.801p 0.53273mV 728043.379p 0.547658mV 728043.837p 0.547658mV 728049.275p 0.545574mV 728063.52p 0.53914mV 728147.16p 0.659658mV 728167.011p 0.632298mV 728216.139p 0.526129mV 728220.017p 0.517193mV 728237.105p 0.451428mV 729015.783p 0.542001mV 729020.508p 0.536054mV 729054.971p 0.478564mV 729074.26p 0.508862mV 730019.806p 0.624951mV 730053.928p 0.726166mV 730073.598p 0.700869mV 730090.487p 0.653862mV 730095.283p 0.644164mV 730100.841p 0.628851mV 730112.642p 0.606172mV 731019.643p 0.560406mV 731024.957p 0.553824mV 731028.297p 0.541006mV 731051.943p 0.570778mV 731052.357p 0.570778mV 731088.954p 0.693951mV 731093.02p 0.715519mV 731094.445p 0.715519mV 732002.755p 0.553171mV 732007.21p 0.552802mV 732032.4p 0.4813mV 733007.853p 0.542781mV 733037.681p 0.583109mV 733043.448p 0.588992mV 733054.074p 0.620314mV 733067.515p 0.679596mV 733071.305p 0.688093mV 733076.999p 0.703653mV 733080.744p 0.726322mV 733085.323p 0.743723mV 734059.97p 0.661197mV 734078.601p 0.702447mV 734083.608p 0.717807mV 735025.131p 0.614543mV 735027.882p 0.614543mV 735033.293p 0.610241mV 735055.449p 0.563068mV 735081.098p 0.374605mV 737025.9p 0.526373mV 737026.048p 0.526373mV 738013.412p 0.593753mV 738037.373p 0.661584mV 738056.201p 0.675866mV 738077.538p 0.677405mV 738094.424p 0.730566mV 738096.051p 0.741878mV 739010.361p 0.583265mV 739016.632p 0.584203mV 739034.465p 0.588342mV 739054.303p 0.597392mV 739098.404p 0.63813mV 739119.043p 0.607257mV 739120.052p 0.597494mV 739132.321p 0.572699mV 739149.65p 0.508535mV 739150.34p 0.487139mV 739164.169p 0.462314mV 739190.62p 0.37363mV 739207.822p 0.351184mV 740035.746p 0.569447mV 740042.447p 0.57593mV 740051.987p 0.595604mV 740120.229p 0.704551mV 741002.058p 0.499344mV 741062.94p 0.327458mV 742000.661p 0.573127mV 742008.52p 0.572145mV 742011.544p 0.577608mV 742018.751p 0.576911mV 742030.985p 0.550612mV 742041.37p 0.531355mV 742055.988p 0.47346mV 743029.135p 0.495226mV 743049.971p 0.472306mV 743058.462p 0.483369mV 743092.561p 0.4942mV 743103.625p 0.511476mV 743122.209p 0.542976mV 743133.476p 0.533065mV 743143.159p 0.522813mV 743159.851p 0.553559mV 743170.402p 0.627917mV 743175.576p 0.657359mV 743178.014p 0.657359mV 743191.071p 0.724177mV 743191.806p 0.724177mV 744029.425p 0.525897mV 744082.706p 0.343421mV 745039.17p 0.650943mV 745063.096p 0.591432mV 745070.441p 0.546864mV 745072.436p 0.546864mV 746000.051p 0.574923mV 746011.667p 0.582632mV 746044.215p 0.559519mV 746045.827p 0.548737mV 746046.678p 0.548737mV 746072.158p 0.513552mV 746109.318p 0.446929mV 746129.73p 0.423853mV 747011.641p 0.531915mV 747052.025p 0.502272mV 747082.302p 0.407269mV 747084.088p 0.407269mV 747098.541p 0.372376mV 748006.01p 0.537077mV 748006.193p 0.537077mV 748035.122p 0.515019mV 748042.796p 0.507724mV 748045.472p 0.493909mV 749002.028p 0.510206mV 749016.827p 0.493483mV 750020.244p 0.502087mV 750037.392p 0.483042mV 750079.005p 0.556013mV 750121.746p 0.580276mV 750152.096p 0.606377mV 750156.079p 0.606518mV 750162.038p 0.613307mV 750163.41p 0.613307mV 750163.622p 0.613307mV 750165.951p 0.626744mV 750188.147p 0.698035mV 750201.31p 0.750421mV 751013.707p 0.573247mV 751014.637p 0.573247mV 751016.265p 0.585229mV 751049.066p 0.630381mV 751049.683p 0.630381mV 751063.997p 0.636106mV 751069.129p 0.639117mV 751084.738p 0.65144mV 751085.355p 0.656669mV 751104.507p 0.713957mV 752037.164p 0.580765mV 752052.108p 0.652345mV 752059.395p 0.67693mV 752067.536p 0.746962mV 753021.575p 0.57932mV 753031.513p 0.588237mV 753036.573p 0.589831mV 753071.815p 0.505189mV 753079.783p 0.494809mV 754004.056p 0.584804mV 754016.217p 0.589445mV 754037.451p 0.565284mV 754078.476p 0.494449mV 754084.448p 0.487982mV 754086.533p 0.487457mV 754144.814p 0.438938mV 754152.069p 0.430855mV 754168.176p 0.460182mV 754182.806p 0.477394mV 754213.736p 0.378841mV 755013.185p 0.530366mV 756010.796p 0.562017mV 756056.707p 0.388206mV 756060.385p 0.367457mV 757021.408p 0.486831mV 757046.634p 0.385744mV 757062.268p 0.330185mV 758009.893p 0.590069mV 758012.151p 0.584086mV 758031.414p 0.54983mV 759037.824p 0.527356mV 759040.169p 0.531453mV 759090.936p 0.754706mV 760005.46p 0.500085mV 760011.664p 0.493475mV 760039.965p 0.461428mV 760057.717p 0.422092mV 760169.27p 0.714945mV 760173.915p 0.748319mV 760174.716p 0.748319mV 761040.153p 0.499814mV 762000.082p 0.549898mV 762004.837p 0.549898mV 762039.609p 0.519931mV 762043.948p 0.501118mV 762046.998p 0.475818mV 763038.884p 0.52409mV 763059.544p 0.472854mV 763059.671p 0.472854mV 763085.038p 0.414316mV 763107.38p 0.402516mV 763140.79p 0.539544mV 763145.379p 0.564413mV 763191.782p 0.758141mV 764024.902p 0.528447mV 764059.005p 0.702875mV 764080.218p 0.748784mV 764084.799p 0.748784mV 765003.72p 0.496443mV 765019.537p 0.516214mV 765069.35p 0.75175mV 766005.799p 0.502235mV 766055.859p 0.546076mV 767000.757p 0.565524mV 767005.565p 0.566495mV 767013.836p 0.573865mV 767052.335p 0.613072mV 767057.603p 0.628539mV 767059.197p 0.628539mV 767078.087p 0.682984mV 767083.229p 0.69524mV 767083.804p 0.69524mV 768011.912p 0.509859mV 768016.738p 0.509265mV 768017.259p 0.509265mV 768067.271p 0.520086mV 768078.5p 0.494446mV 768102.964p 0.452646mV 768107.083p 0.458972mV 768107.715p 0.458972mV 768164.637p 0.510003mV 768184.808p 0.641671mV 768199.571p 0.733791mV 769001.427p 0.514213mV 769014.394p 0.519598mV 769024.545p 0.536704mV 769029.62p 0.548195mV 769052.996p 0.573813mV 769061.302p 0.565646mV 769102.306p 0.5104mV 769117.043p 0.449934mV 769136.965p 0.336476mV 770026.594p 0.517937mV 770037.285p 0.533978mV 770058.796p 0.589727mV 771038.253p 0.691789mV 771044.553p 0.713945mV 771046.45p 0.743227mV 772061.67p 0.449028mV 772088.558p 0.418949mV 773002.887p 0.56879mV 773003.39p 0.56879mV 773014.038p 0.563041mV 773021.091p 0.557733mV 773025.622p 0.545753mV 773028.164p 0.545753mV 773056.457p 0.49087mV 773074.176p 0.487665mV 773125.505p 0.38692mV 774029.769p 0.601802mV 774047.302p 0.630647mV 774064.707p 0.600534mV 774092.326p 0.441054mV 774100.378p 0.365261mV 775002.94p 0.549368mV 775038.16p 0.549231mV 775041.736p 0.541905mV 775047.511p 0.540876mV 775067.289p 0.574189mV 775080.652p 0.647262mV 775086.598p 0.67227mV 775087.62p 0.67227mV 775096.541p 0.70547mV 775116.535p 0.720617mV 775123.971p 0.720765mV 775128.534p 0.728194mV 775138.664p 0.752527mV 776011.846p 0.607702mV 776028.842p 0.614827mV 776029.415p 0.614827mV 776069.104p 0.608221mV 776088.094p 0.650871mV 777020.498p 0.586142mV 777087.136p 0.553628mV 778038.927p 0.585447mV 778060.187p 0.597653mV 778071.453p 0.633315mV 778103.831p 0.702584mV 778110.37p 0.748503mV 779004.358p 0.588624mV 779054.047p 0.756637mV 779054.069p 0.756637mV 780004.358p 0.550992mV 780015.371p 0.547795mV 780020.199p 0.542519mV 780020.658p 0.542519mV 780043.665p 0.508217mV 780049.284p 0.496079mV 780076.654p 0.42065mV 780079.037p 0.42065mV 780087.338p 0.419253mV 780128.608p 0.326953mV 781004.882p 0.601821mV 781031.164p 0.673038mV 781038.752p 0.700256mV 782001.796p 0.529163mV 782013.264p 0.533966mV 782036.867p 0.515658mV 783018.58p 0.585671mV 783036.638p 0.591649mV 783047.014p 0.577315mV 783053.803p 0.56107mV 783061.03p 0.510093mV 783077.916p 0.448382mV 785035.317p 0.405463mV 785049.538p 0.352094mV 786021.83p 0.602499mV 786042.906p 0.585188mV 786061.293p 0.635224mV 786075.14p 0.7304mV 787002.84p 0.553452mV 787021.097p 0.592905mV 787068.561p 0.703682mV 787075.328p 0.76025mV 788082.365p 0.729351mV 788086.971p 0.770597mV 788087.942p 0.770597mV 789000.527p 0.598319mV 789016.335p 0.591674mV 789016.769p 0.591674mV 789035.81p 0.582587mV 789044.054p 0.577897mV 789173.353p 0.539107mV 789189.019p 0.631048mV 789199.223p 0.695709mV 790001.444p 0.499165mV 790007.202p 0.498415mV 790058.841p 0.453658mV 791080.606p 0.40765mV 792027.27p 0.552402mV 792126.899p 0.417288mV 792142.187p 0.388531mV 792154.698p 0.341886mV 793013.262p 0.495297mV 793020.56p 0.473915mV 794006.016p 0.563419mV 794009.098p 0.563419mV 794012.065p 0.558038mV 794020.903p 0.553799mV 794025.37p 0.554912mV 794038.355p 0.563519mV 794054.326p 0.580163mV 794074.226p 0.676298mV 795015.457p 0.512356mV 796033.573p 0.634584mV 796048.115p 0.623374mV 796054.514p 0.608141mV 796093.102p 0.548042mV 796116.681p 0.513687mV 796168.024p 0.496864mV 796182.062p 0.526048mV 796204.068p 0.541353mV 796208.031p 0.541922mV 796238.808p 0.525682mV 796262.363p 0.531722mV 796279.828p 0.51083mV 796330.246p 0.616521mV 796330.722p 0.616521mV 796332.982p 0.616521mV 796339.935p 0.640312mV 796341.856p 0.670808mV 797001.034p 0.496607mV 797042.4p 0.593697mV 797093.945p 0.501976mV 797162.317p 0.439899mV 797209.724p 0.674761mV 797220.222p 0.771684mV 798011.842p 0.597615mV 798044.693p 0.525085mV 798047.471p 0.501626mV 798050.674p 0.47171mV 798056.455p 0.447787mV 798060.599p 0.429656mV 799001.524p 0.548637mV 799030.717p 0.581458mV 799048.04p 0.589784mV 799076.228p 0.504595mV 799096.896p 0.445319mV 800002.239p 0.603543mV 800043.818p 0.634355mV 801010.221p 0.580029mV 801030.924p 0.609025mV 801050.522p 0.668695mV 801052.8p 0.668695mV 801054.096p 0.668695mV 801056.357p 0.697482mV 802006.779p 0.517403mV 802091.554p 0.350411mV 803002.208p 0.584585mV 803012.651p 0.589568mV 803031.292p 0.551894mV 804000.496p 0.532825mV 804048.891p 0.639521mV 804075.987p 0.758576mV 804076.444p 0.758576mV 806051.413p 0.557112mV 806081.593p 0.698908mV 807030.708p 0.609105mV 807041.891p 0.667931mV 807056.438p 0.732544mV 807059.772p 0.732544mV 807068.757p 0.761823mV 808010.543p 0.559874mV 808014.491p 0.559874mV 808034.663p 0.545476mV 808037.01p 0.545099mV 808051.65p 0.543745mV 808064.139p 0.536231mV 809049.086p 0.5238mV 809089.612p 0.454033mV 809122.005p 0.43695mV 809142.527p 0.452507mV 809166.263p 0.455286mV 809170.112p 0.445279mV 809174.68p 0.445279mV 809192.066p 0.411324mV 810082.338p 0.65301mV 810086.526p 0.667082mV 810087.786p 0.667082mV 811023.183p 0.486138mV 811090.28p 0.70688mV 811095.904p 0.742481mV 812006.384p 0.523096mV 812006.768p 0.523096mV 812044.122p 0.510719mV 812095.08p 0.554785mV 812099.845p 0.554785mV 812101.413p 0.557503mV 812143.495p 0.660523mV 812158.317p 0.716132mV 813075.341p 0.527298mV 813103.863p 0.581228mV 813123.054p 0.533144mV 813141.151p 0.421823mV 813141.258p 0.421823mV 814002.174p 0.526851mV 814049.526p 0.43005mV 814075.665p 0.330151mV 815022.294p 0.499556mV 815023.092p 0.499556mV 815142.691p 0.327145mV 816035.009p 0.57361mV 816040.51p 0.580366mV 816041.53p 0.580366mV 816042.011p 0.580366mV 816042.109p 0.580366mV 816065.537p 0.547362mV 816096.394p 0.369399mV 817010.679p 0.493301mV 817021.327p 0.461853mV 817127.605p 0.610535mV 817152.501p 0.636055mV 817158.869p 0.631335mV 817178.454p 0.642916mV 817188.93p 0.633324mV 817196.391p 0.625904mV 817201.992p 0.632361mV 817218.422p 0.642156mV 817221.563p 0.650696mV 817263.005p 0.721088mV 817264.345p 0.721088mV 818019.056p 0.561691mV 818042.814p 0.408383mV 818047.044p 0.357834mV 819064.533p 0.453713mV 820004.065p 0.523953mV 820008.452p 0.524635mV 820009.633p 0.524635mV 820013.587p 0.531453mV 820030.459p 0.49435mV 820042.162p 0.461986mV 820053.505p 0.415272mV 820064.97p 0.390775mV 820084.388p 0.367696mV 821011.191p 0.555587mV 821050.136p 0.427538mV 822014.349p 0.551491mV 822017.104p 0.564002mV 822020.386p 0.582824mV 822028.286p 0.608035mV 822050.368p 0.695766mV 822067.154p 0.764497mV 823018.477p 0.569493mV 823022.77p 0.588971mV 824081.444p 0.734221mV 825004.828p 0.556248mV 825009.657p 0.555859mV 825025.146p 0.516666mV 825025.212p 0.516666mV 825079.568p 0.491191mV 825080.596p 0.4812mV 825082.606p 0.4812mV 825142.857p 0.514693mV 825144.425p 0.514693mV 825171.931p 0.664704mV 825197.476p 0.730623mV 825200.559p 0.745439mV 826002.715p 0.579302mV 826007.988p 0.578278mV 826023.402p 0.601528mV 826028.374p 0.601372mV 827005.705p 0.560416mV 827017.716p 0.56657mV 827019.931p 0.56657mV 827031.538p 0.554435mV 827034.731p 0.554435mV 827053.003p 0.49244mV 828004.86p 0.522043mV 828035.777p 0.568689mV 828036.123p 0.568689mV 828056.14p 0.61358mV 828072.726p 0.612527mV 828086.407p 0.583713mV 828089.497p 0.583713mV 828093.615p 0.56634mV 828103.835p 0.55102mV 828117.711p 0.575591mV 828167.759p 0.68139mV 829015.085p 0.584107mV 829030.727p 0.558228mV 829101.859p 0.647864mV 829102.74p 0.647864mV 829115.662p 0.761624mV 830041.043p 0.49694mV 830042.191p 0.49694mV 830062.978p 0.489394mV 830068.435p 0.486552mV 832003.914p 0.513583mV 832059.166p 0.561062mV 832081.104p 0.624893mV 832097.274p 0.619691mV 832108.497p 0.641523mV 832130.245p 0.740614mV 833027.673p 0.640138mV 833028.128p 0.640138mV 833033.906p 0.660949mV 835037.014p 0.632116mV 835041.39p 0.628268mV 835082.732p 0.744299mV 836004.662p 0.582447mV 836034.286p 0.562791mV 836040.716p 0.544723mV 836041.249p 0.544723mV 836062.972p 0.457811mV 836076.915p 0.373137mV 837020.588p 0.533149mV 837031.768p 0.540448mV 837049.705p 0.522395mV 837083.467p 0.351965mV 838023.904p 0.569536mV 838029.728p 0.568978mV 838038.36p 0.574528mV 838066.31p 0.556005mV 838066.372p 0.556005mV 838097.793p 0.423948mV 840008.381p 0.577484mV 840027.655p 0.593917mV 840031.343p 0.589167mV 840032.365p 0.589167mV 840048.34p 0.538642mV 840064.386p 0.494932mV 840066.038p 0.484178mV 841007.948p 0.565642mV 841011.68p 0.571355mV 842011.485p 0.590157mV 842014.564p 0.590157mV 842042.19p 0.502941mV 842064.313p 0.429248mV 843000.962p 0.575101mV 843014.032p 0.58255mV 843027.458p 0.617193mV 843055.768p 0.691744mV 843059.403p 0.691744mV 843066.27p 0.709972mV 843099.7p 0.739667mV 844028.909p 0.575982mV 844036.5p 0.607888mV 844038.015p 0.607888mV 844048.732p 0.615706mV 844061.774p 0.633634mV 844065.768p 0.648908mV 844075.518p 0.687414mV 845034.133p 0.628014mV 845034.502p 0.628014mV 845040.283p 0.640778mV 845068.572p 0.718024mV 845075.118p 0.716605mV 845111.631p 0.760401mV 846020.371p 0.54629mV 846038.999p 0.528338mV 846039.351p 0.528338mV 846045.751p 0.484565mV 846079.335p 0.431286mV 846113.174p 0.386874mV 846153.838p 0.442136mV 846158.372p 0.437732mV 846174.804p 0.457958mV 846179.642p 0.475874mV 846181.575p 0.486936mV 846192.968p 0.51401mV 846206.343p 0.543071mV 846210.142p 0.565002mV 846248.485p 0.710789mV 846254.313p 0.73556mV 846255.335p 0.767555mV 847001.675p 0.550625mV 847037.395p 0.61153mV 847063.813p 0.728983mV 847071.483p 0.770676mV 847074.117p 0.770676mV 848032.895p 0.494317mV 849015.243p 0.553996mV 849025.363p 0.584185mV 849028.605p 0.584185mV 849036.948p 0.627491mV 849072.128p 0.717034mV 849076.66p 0.734868mV 849078.676p 0.734868mV 849079.433p 0.734868mV 850015.512p 0.552249mV 850024.064p 0.558814mV 850045.671p 0.687767mV 851012.049p 0.604036mV 851042.284p 0.581559mV 851071.168p 0.528171mV 851139.228p 0.496871mV 851173.725p 0.425472mV 851184.097p 0.374045mV 852001.509p 0.547603mV 852035.952p 0.545714mV 852069.592p 0.632414mV 852080.148p 0.651743mV 852091.6p 0.665443mV 852103.69p 0.669306mV 852122.695p 0.648335mV 852139.208p 0.620921mV 852139.234p 0.620921mV 852152.406p 0.554208mV 852156.835p 0.528281mV 852184.269p 0.45298mV 852185.618p 0.437914mV 852206.266p 0.370441mV 853027.123p 0.508796mV 854007.431p 0.583442mV 854037.46p 0.690073mV 854043.329p 0.723212mV 854048.373p 0.763463mV 855035.105p 0.619495mV 855054.072p 0.649764mV 855064.366p 0.64965mV 855084.609p 0.669718mV 855113.443p 0.728691mV 855125.23p 0.774239mV 856011.741p 0.512401mV 856018.561p 0.524533mV 856035.917p 0.558955mV 856036.574p 0.558955mV 856047.859p 0.563661mV 856048.84p 0.563661mV 856053.221p 0.556681mV 856060.396p 0.549236mV 856066.644p 0.548725mV 856070.385p 0.55451mV 856110.313p 0.681357mV 856114.957p 0.681357mV 856119.675p 0.696094mV 856133.314p 0.720599mV 856146.249p 0.723138mV 856146.35p 0.723138mV 856164.317p 0.692059mV 856207.473p 0.671415mV 856215.565p 0.692487mV 856248.77p 0.676694mV 856262.102p 0.671245mV 856273.178p 0.648557mV 856274.715p 0.648557mV 856291.814p 0.585775mV 856297.785p 0.567942mV 856311.168p 0.47751mV 856324.168p 0.422624mV 857017.113p 0.534862mV 857035.141p 0.592533mV 857037.509p 0.592533mV 857046.688p 0.659571mV 858022.844p 0.574872mV 858025.944p 0.574634mV 858033.576p 0.568254mV 858051.836p 0.581888mV 858098.799p 0.689531mV 859009.783p 0.496852mV 859014.66p 0.502476mV 859072.343p 0.553846mV 859108.849p 0.681967mV 859109.425p 0.681967mV 859125.348p 0.76065mV 860023.136p 0.551338mV 861008.793p 0.558209mV 861078.237p 0.414746mV 862036.907p 0.667352mV 863015.054p 0.567069mV 863015.827p 0.567069mV 863038.489p 0.528114mV 863040.644p 0.521516mV 863047.03p 0.508481mV 863048.008p 0.508481mV 864000.675p 0.514291mV 864037.975p 0.375362mV 865040.571p 0.568191mV 865068.538p 0.56685mV 865071.814p 0.563309mV 865073.007p 0.563309mV 865084.863p 0.537621mV 865092.363p 0.524587mV 865106.279p 0.513492mV 865108.421p 0.513492mV 866000.5p 0.59427mV 866014.311p 0.588975mV 866025.405p 0.586185mV 866027.818p 0.586185mV 867028.554p 0.573555mV 867059.547p 0.638344mV 867079.636p 0.602613mV 867103.904p 0.636341mV 867108.866p 0.643048mV 867117.882p 0.639303mV 867164.638p 0.627749mV 867172.425p 0.623169mV 867173.676p 0.623169mV 867174.862p 0.623169mV 867175.013p 0.612194mV 867181.184p 0.607965mV 867193.467p 0.619526mV 867199.008p 0.635306mV 867224.3p 0.766898mV 868046.499p 0.577829mV 868064.417p 0.640637mV 868070.933p 0.699133mV 869009.372p 0.569953mV 869076.693p 0.652756mV 869082.15p 0.640468mV 869097.571p 0.582057mV 869107.081p 0.542825mV 869120.461p 0.493619mV 870001.448p 0.602463mV 870036.95p 0.537417mV 870084.708p 0.525127mV 870111.308p 0.58027mV 870125.332p 0.599553mV 870127.036p 0.599553mV 870162.823p 0.62451mV 870178.422p 0.642293mV 870198.215p 0.703237mV 870200.686p 0.717233mV 870205.047p 0.738419mV 870212.943p 0.754435mV 871062.735p 0.531724mV 871084.363p 0.609701mV 871091.987p 0.649434mV 871103.117p 0.703742mV 871112.22p 0.761158mV 872028.114p 0.565073mV 872046.339p 0.639367mV 872128.181p 0.670897mV 872156.344p 0.677263mV 872163.039p 0.661582mV 872195.655p 0.504225mV 872207.401p 0.458748mV 872216.501p 0.411515mV 872222.298p 0.396272mV 872229.612p 0.373918mV 873011.404p 0.545434mV 873011.607p 0.545434mV 873021.097p 0.525222mV 873030.933p 0.529804mV 873051.271p 0.537259mV 873052.612p 0.537259mV 873055.088p 0.548287mV 873077.206p 0.592175mV 873084.211p 0.609714mV 873124.35p 0.703598mV 873137.962p 0.724877mV 873138.56p 0.724877mV 873146.44p 0.758724mV 874062.038p 0.460764mV 874066.601p 0.4671mV 874067.953p 0.4671mV 875029.819p 0.604289mV 875031.796p 0.610529mV 875047.741p 0.656672mV 877009.227p 0.597321mV 877019.554p 0.591883mV 877034.574p 0.595237mV 877035.486p 0.584376mV 877039.235p 0.584376mV 877062.967p 0.514291mV 877077.763p 0.489413mV 877091.294p 0.480495mV 877092.405p 0.480495mV 877094.546p 0.480495mV 877095.002p 0.468332mV 877102.581p 0.462018mV 877104.645p 0.462018mV 877110.6p 0.441525mV 877125.194p 0.402793mV 877128.493p 0.402793mV 878012.468p 0.526334mV 878076.184p 0.489932mV 878095.807p 0.474595mV 878102.489p 0.475942mV 878111.246p 0.496073mV 878149.279p 0.541999mV 879012.673p 0.504275mV 881016.526p 0.521523mV 881037.339p 0.478903mV 881038.911p 0.478903mV 882036.001p 0.51287mV 882038.729p 0.51287mV 882073.605p 0.563641mV 882103.022p 0.675941mV 882115.272p 0.767266mV 882116.064p 0.767266mV 882117.882p 0.767266mV 883033.31p 0.580356mV 883094.066p 0.609308mV 883097.531p 0.614852mV 883106.331p 0.645966mV 883110.003p 0.659072mV 883113.837p 0.659072mV 883129.598p 0.714917mV 883131.898p 0.731038mV 884003.929p 0.541787mV 884026.743p 0.53704mV 884066.752p 0.512374mV 885015.684p 0.562641mV 885019.832p 0.562641mV 885040.825p 0.617156mV 885044.763p 0.617156mV 886003.207p 0.52035mV 886012.073p 0.525845mV 886013.333p 0.525845mV 886035.854p 0.558851mV 886050.888p 0.59331mV 886071.733p 0.604344mV 886126.183p 0.394666mV 887034.499p 0.56691mV 887046.901p 0.623568mV 887049.99p 0.623568mV 887062.097p 0.702335mV 888000.408p 0.50678mV 888033.794p 0.594121mV 889003.859p 0.553409mV 889012.442p 0.559999mV 889014.344p 0.559999mV 889021.381p 0.579322mV 889036.316p 0.612615mV 889055.766p 0.657894mV 889062.227p 0.655007mV 889085.804p 0.656544mV 889090.92p 0.657465mV 889109.798p 0.639175mV 889131.307p 0.637275mV 889160.12p 0.729016mV 889169.677p 0.733913mV 889193.742p 0.74528mV 889208.899p 0.730013mV 889216.562p 0.731712mV 889216.571p 0.731712mV 889219.784p 0.731712mV 889224.808p 0.731133mV 889234.623p 0.751986mV 889238.722p 0.773447mV 890019.753p 0.603094mV 890021.372p 0.610178mV 890115.332p 0.703613mV 890167.737p 0.49272mV 891027.033p 0.586159mV 891030.515p 0.581606mV 891033.246p 0.581606mV 891042.38p 0.592049mV 891044.184p 0.592049mV 891067.816p 0.556213mV 891076.815p 0.556936mV 891080.641p 0.566791mV 891124.633p 0.483737mV 891134.254p 0.458235mV 891157.113p 0.348984mV 891176.933p 0.343677mV 891178.117p 0.343677mV 891194.274p 0.341352mV 891200.331p 0.347746mV 892056.681p 0.524469mV 892075.003p 0.542757mV 893001.265p 0.570545mV 893038.436p 0.53607mV 893041.091p 0.541984mV 893041.679p 0.541984mV 893062.485p 0.590456mV 893077.894p 0.609325mV 893090.166p 0.63768mV 893096.849p 0.63966mV 893096.931p 0.63966mV 893101.537p 0.635915mV 893124.009p 0.651588mV 894020.831p 0.509058mV 894023.146p 0.509058mV 894040.904p 0.502699mV 894050.068p 0.529175mV 894063.154p 0.579946mV 894064.971p 0.579946mV 894066.337p 0.602124mV 895013.214p 0.54023mV 895028.158p 0.483634mV 896055.507p 0.404579mV 897029.441p 0.458994mV 898030.138p 0.550986mV 898031.499p 0.550986mV 898062.743p 0.531794mV 898063.192p 0.531794mV 898091.785p 0.421203mV 899002.496p 0.556768mV 899003.969p 0.556768mV 899033.947p 0.572104mV 899062.524p 0.503668mV 900011.974p 0.510384mV 900013.102p 0.510384mV 900017.956p 0.497946mV 900019.042p 0.497946mV 900048.308p 0.473236mV 901011.735p 0.553891mV 901020.932p 0.52296mV 901026.489p 0.510604mV 901037.965p 0.466409mV 902003.85p 0.593206mV 902053.732p 0.475058mV 902078.094p 0.343636mV 903046.585p 0.645154mV 903048.364p 0.645154mV 903049.764p 0.645154mV 903054.535p 0.6645mV 903068.37p 0.688981mV 903083.97p 0.677231mV 903103.364p 0.74404mV 904065.388p 0.630453mV 904092.392p 0.737767mV 904095.391p 0.755522mV 905026.765p 0.534817mV 905033.824p 0.541055mV 905043.936p 0.534379mV 905060.13p 0.570535mV 905070.472p 0.588526mV 905070.771p 0.588526mV 905075.586p 0.60094mV 905113.707p 0.621697mV 905116.343p 0.624572mV 905123.336p 0.634184mV 905130.063p 0.63603mV 905147.063p 0.646047mV 905152.029p 0.658883mV 905153.544p 0.658883mV 906000.389p 0.567115mV 906004.858p 0.567115mV 906013.618p 0.575397mV 906026.72p 0.560461mV 906055.706p 0.514096mV 906073.122p 0.480242mV 906074.926p 0.480242mV 906082.735p 0.462121mV 906095.836p 0.465624mV 906108.975p 0.454808mV 906143.375p 0.446214mV 906156.698p 0.40397mV 906168.404p 0.340695mV 907009.63p 0.557193mV 907023.449p 0.585079mV 907023.894p 0.585079mV 907024.033p 0.585079mV 907062.864p 0.600632mV 907071.443p 0.613637mV 907090.164p 0.669598mV 907092.791p 0.669598mV 907104.679p 0.676181mV 907116.962p 0.65751mV 907120.453p 0.64858mV 907133.358p 0.613889mV 908001.07p 0.555492mV 908013.39p 0.549924mV 908027.644p 0.5196mV 908057.199p 0.536704mV 908075.64p 0.583119mV 908094.34p 0.619296mV 908098.902p 0.632032mV 908111.84p 0.647996mV 908112.979p 0.647996mV 908118.518p 0.662798mV 908121.673p 0.671944mV 908128.6p 0.688061mV 909011.346p 0.532058mV 909032.713p 0.559782mV 909036.83p 0.5603mV 909056.386p 0.562901mV 909073.12p 0.565539mV 909114.754p 0.381688mV 910017.176p 0.598308mV 910049.403p 0.628785mV 910052.324p 0.638268mV 911001.593p 0.571857mV 911010.28p 0.564777mV 911096.838p 0.436835mV 911103.208p 0.459476mV 911117.327p 0.498611mV 911138.89p 0.579256mV 911157.603p 0.585149mV 911177.498p 0.645214mV 911188.649p 0.684078mV 911222.165p 0.712177mV 911258.006p 0.746836mV 911270.081p 0.733938mV 911276.521p 0.732087mV 911316.548p 0.680788mV 911365.375p 0.680507mV 911365.937p 0.680507mV 911369.556p 0.680507mV 911396.072p 0.625075mV 911396.234p 0.625075mV 911402.006p 0.613033mV 911413.119p 0.60915mV 911422.367p 0.619347mV 911426.102p 0.628198mV 911430.197p 0.643772mV 911468.346p 0.631574mV 911482.766p 0.575258mV 911495.265p 0.527691mV 911507.876p 0.527313mV 911527.001p 0.600642mV 911531.757p 0.634799mV 912008.444p 0.535185mV 912047.778p 0.539749mV 912109.137p 0.372321mV 913035.069p 0.641312mV 913039.871p 0.641312mV 913041.532p 0.663432mV 913058.897p 0.721194mV 913060.172p 0.746336mV 913063.032p 0.746336mV 914005.45p 0.589043mV 914005.776p 0.589043mV 914005.952p 0.589043mV 914008.333p 0.589043mV 914022.905p 0.630245mV 914048.037p 0.695818mV 914053.077p 0.695007mV 914081.342p 0.614492mV 915000.148p 0.539193mV 915014.862p 0.547047mV 915026.546p 0.580619mV 916009.301p 0.562983mV 916024.407p 0.537585mV 917008.169p 0.564887mV 917047.873p 0.561648mV 917107.787p 0.381584mV 917122.142p 0.385396mV 918013.261p 0.545609mV 918025.91p 0.586946mV 918031.001p 0.605104mV 918040.99p 0.63593mV 918044.105p 0.63593mV 919003.434p 0.507927mV 919009.893p 0.507305mV 919016.009p 0.486371mV 919035.899p 0.414647mV 919057.275p 0.33137mV 919059.29p 0.33137mV 920031.945p 0.434201mV 920034.356p 0.434201mV 921001.622p 0.586319mV 921004.319p 0.586319mV 921019.15p 0.571011mV 921019.713p 0.571011mV 921032.332p 0.500608mV 921034.602p 0.500608mV 922000.788p 0.597994mV 922002.196p 0.597994mV 922004.468p 0.597994mV 922016.431p 0.615276mV 922025.533p 0.659937mV 922033.039p 0.679864mV 923006.457p 0.576537mV 924042.72p 0.354004mV 924044.357p 0.354004mV 925010.898p 0.556203mV 925097.947p 0.525652mV 926004.82p 0.514448mV 926033.072p 0.467046mV 926066.483p 0.435258mV 926099.131p 0.467865mV 926168.767p 0.379795mV 927013.97p 0.586309mV 927026.436p 0.556197mV 927057.569p 0.426139mV 927073.65p 0.382103mV 929011.078p 0.562874mV 929054.179p 0.733447mV 930009.707p 0.543449mV 930028.525p 0.606357mV 930046.949p 0.698416mV 930052.583p 0.707516mV 930052.851p 0.707516mV 930067.343p 0.728127mV 930067.432p 0.728127mV 931003.055p 0.528806mV 931017.702p 0.536321mV 931099.502p 0.431419mV 931130.793p 0.353289mV 932002.358p 0.561995mV 932007.898p 0.561383mV 932010.761p 0.554546mV 932050.263p 0.419378mV 933013.114p 0.494033mV 933018.717p 0.481644mV 933020.649p 0.46261mV 933045.496p 0.339017mV 934012.57p 0.503003mV 934024.571p 0.483355mV 934044.989p 0.464551mV 935002.0p 0.569025mV 935028.585p 0.555073mV 935041.767p 0.517629mV 935042.426p 0.517629mV 935067.564p 0.46405mV 935083.462p 0.456988mV 936004.892p 0.567483mV 936041.18p 0.564107mV 936061.954p 0.608453mV 936062.383p 0.608453mV 936063.815p 0.608453mV 936077.113p 0.622587mV 936088.016p 0.636195mV 936091.456p 0.634323mV 936112.182p 0.670028mV 936116.515p 0.677386mV 936119.053p 0.677386mV 936139.097p 0.652119mV 936163.395p 0.595018mV 936163.898p 0.595018mV 936193.3p 0.587545mV 936197.491p 0.590527mV 936214.083p 0.600928mV 936252.075p 0.618163mV 936253.357p 0.618163mV 936269.902p 0.65974mV 936271.899p 0.674626mV 936293.778p 0.679272mV 936311.752p 0.672251mV 936314.533p 0.672251mV 936340.662p 0.709788mV 936357.607p 0.743168mV 936379.096p 0.733581mV 936421.708p 0.725622mV 936481.682p 0.732974mV 936482.606p 0.732974mV 936485.058p 0.758851mV 937039.779p 0.517535mV 937074.866p 0.460463mV 937076.83p 0.457898mV 937077.661p 0.457898mV 937081.475p 0.448493mV 938016.94p 0.532927mV 938034.748p 0.481358mV 938079.039p 0.359678mV 938080.414p 0.345088mV 938098.954p 0.33092mV 938112.228p 0.347704mV 938147.335p 0.352015mV 938153.834p 0.356487mV 939000.678p 0.598318mV 939007.805p 0.597387mV 940015.565p 0.616584mV 940026.977p 0.661332mV 940033.073p 0.693875mV 940040.749p 0.742479mV 940049.534p 0.771389mV 941011.124p 0.586423mV 941028.519p 0.572612mV 941036.054p 0.570741mV 941060.163p 0.641423mV 941074.358p 0.693614mV 941084.265p 0.748777mV 941084.557p 0.748777mV 941084.9p 0.748777mV 942000.315p 0.517244mV 942012.854p 0.522356mV 942038.589p 0.579214mV 942072.28p 0.768986mV 943008.346p 0.542696mV 943021.505p 0.526898mV 943031.417p 0.492767mV 943031.485p 0.492767mV 943047.965p 0.442631mV 944015.25p 0.502821mV 944020.557p 0.483559mV 944030.124p 0.425149mV 945000.511p 0.563667mV 945022.258p 0.603704mV 946006.939p 0.560491mV 946027.145p 0.558807mV 946036.99p 0.577324mV 946053.835p 0.653347mV 946070.348p 0.749494mV 947012.389p 0.610527mV 947043.691p 0.691728mV 947131.779p 0.695298mV 947132.789p 0.695298mV 947133.251p 0.695298mV 947140.17p 0.737151mV 947141.708p 0.737151mV 948026.583p 0.624462mV 948049.309p 0.707112mV 948049.33p 0.707112mV 948059.866p 0.746891mV 949016.852p 0.603907mV 949030.188p 0.633473mV 949069.476p 0.730946mV 950022.064p 0.53392mV 950030.696p 0.502958mV 950048.147p 0.470605mV 950070.172p 0.377399mV 951001.405p 0.57914mV 951014.071p 0.586286mV 951020.349p 0.594215mV 951038.37p 0.592253mV 951064.183p 0.522515mV 951090.837p 0.414781mV 951104.958p 0.370512mV 951106.584p 0.356298mV 952003.954p 0.553032mV 952044.997p 0.639788mV 952055.637p 0.687944mV 952057.601p 0.687944mV 952074.515p 0.711664mV 952078.276p 0.717265mV 952097.614p 0.700263mV 952132.392p 0.65798mV 952137.063p 0.649908mV 952179.5p 0.604066mV 952184.31p 0.606278mV 952187.792p 0.602539mV 952197.441p 0.577224mV 952281.238p 0.382mV 952288.729p 0.391739mV 952304.7p 0.377514mV 953017.177p 0.550792mV 954004.378p 0.58861mV 954023.313p 0.617605mV 954048.089p 0.567611mV 954056.608p 0.543525mV 954085.039p 0.430777mV 954091.069p 0.426014mV 954100.733p 0.407948mV 954111.255p 0.374031mV 955007.068p 0.536957mV 955009.21p 0.536957mV 955012.862p 0.543394mV 955029.278p 0.524525mV 955032.046p 0.518113mV 955054.184p 0.465141mV 955064.833p 0.430149mV 955069.27p 0.402355mV 956055.207p 0.581642mV 956064.414p 0.576388mV 956101.945p 0.566643mV 956109.407p 0.569428mV 956116.074p 0.556427mV 957004.325p 0.558509mV 957012.019p 0.566511mV 957021.597p 0.599994mV 958012.096p 0.523086mV 958018.21p 0.522955mV 958037.901p 0.533436mV 958090.319p 0.689867mV 958092.863p 0.689867mV 958099.182p 0.703808mV 958122.633p 0.756767mV 958124.104p 0.756767mV 958124.922p 0.756767mV 959003.835p 0.506763mV 959118.101p 0.665108mV 959130.503p 0.68847mV 959133.749p 0.68847mV 959133.997p 0.68847mV 959145.963p 0.750495mV 960010.722p 0.584807mV 960020.747p 0.590804mV 960028.186p 0.603578mV 960043.596p 0.60596mV 960074.556p 0.524514mV 960105.648p 0.518324mV 960119.86p 0.513813mV 960193.835p 0.633457mV 960194.926p 0.633457mV 960231.096p 0.683487mV 960232.885p 0.683487mV 960238.239p 0.717187mV 960239.792p 0.717187mV 960243.788p 0.745469mV 961045.552p 0.544154mV 961068.67p 0.662954mV 961073.689p 0.693429mV 961082.629p 0.762963mV 962000.617p 0.549799mV 962006.807p 0.549836mV 962013.152p 0.556174mV 962018.56p 0.556209mV 962019.327p 0.556209mV 962024.481p 0.562584mV 962038.132p 0.582065mV 962043.685p 0.601361mV 962044.652p 0.601361mV 962067.062p 0.684696mV 962100.858p 0.703812mV 962111.784p 0.693771mV 962115.423p 0.6933mV 962129.675p 0.688829mV 962161.229p 0.570522mV 962168.103p 0.539618mV 962174.094p 0.502541mV 962190.321p 0.326052mV 964003.072p 0.579679mV 964036.354p 0.627272mV 964038.42p 0.627272mV 964047.246p 0.650529mV 964048.408p 0.650529mV 964048.844p 0.650529mV 964078.268p 0.749775mV 964079.645p 0.749775mV 964080.258p 0.752341mV 964091.301p 0.767419mV 965002.602p 0.516252mV 965002.671p 0.516252mV 965031.29p 0.54775mV 965050.527p 0.595523mV 965062.975p 0.626534mV 965064.363p 0.626534mV 965068.716p 0.639403mV 965101.367p 0.774533mV 966062.216p 0.459424mV 966078.028p 0.406367mV 967024.19p 0.56512mV 967047.021p 0.560975mV 967056.819p 0.545708mV 967096.044p 0.483709mV 968013.913p 0.513833mV 968028.629p 0.464909mV 968032.224p 0.443681mV 968033.061p 0.443681mV 969039.003p 0.594773mV 969065.449p 0.742849mV 970000.129p 0.595962mV 970013.143p 0.590636mV 970028.468p 0.550029mV 970046.477p 0.530524mV 970056.211p 0.526782mV 970057.008p 0.526782mV 970066.701p 0.547663mV 970077.212p 0.568183mV 970085.88p 0.601468mV 970099.271p 0.635668mV 970133.925p 0.764391mV 971010.498p 0.519492mV 971032.831p 0.541361mV 971042.093p 0.54523mV 971048.3p 0.556528mV 971068.018p 0.627448mV 971076.637p 0.658295mV 971079.808p 0.658295mV 971090.29p 0.699875mV 972020.997p 0.516759mV 972023.157p 0.516759mV 972043.927p 0.375273mV 973025.955p 0.598089mV 973033.217p 0.62915mV 974021.806p 0.536386mV 974032.439p 0.506269mV 974081.43p 0.381714mV 975010.566p 0.535837mV 975015.742p 0.523614mV 975015.874p 0.523614mV 975017.489p 0.523614mV 975024.976p 0.517604mV 975025.63p 0.505127mV 975046.524p 0.515545mV 975060.39p 0.548831mV 975063.564p 0.548831mV 976027.377p 0.550785mV 976028.095p 0.550785mV 977020.579p 0.539462mV 977027.337p 0.526681mV 978003.987p 0.567714mV 978004.403p 0.567714mV 978015.51p 0.550482mV 978019.826p 0.550482mV 978039.291p 0.490306mV 979048.555p 0.5675mV 980009.684p 0.569963mV 980026.38p 0.632131mV 981032.843p 0.488684mV 981039.803p 0.47371mV 982002.103p 0.552903mV 982026.856p 0.53558mV 982055.558p 0.368719mV 983078.92p 0.470869mV 984020.967p 0.516102mV 984031.895p 0.49456mV 984073.735p 0.442331mV 984077.762p 0.448834mV 985006.233p 0.535907mV 985024.732p 0.532571mV 985037.321p 0.534415mV 985038.279p 0.534415mV 985089.823p 0.740888mV 986008.449p 0.502291mV 986009.804p 0.502291mV 986032.174p 0.558385mV 986075.609p 0.727927mV 987011.781p 0.572357mV 987043.008p 0.576921mV 987068.041p 0.591991mV 987076.767p 0.575677mV 987124.0p 0.402349mV 988001.09p 0.537081mV 988022.781p 0.509163mV 988037.353p 0.44847mV 989008.382p 0.600205mV 989010.176p 0.606134mV 989027.21p 0.625926mV 989031.729p 0.645853mV 990004.477p 0.541394mV 990039.319p 0.609368mV 990086.674p 0.685299mV 990089.547p 0.685299mV 990098.924p 0.669981mV 990101.901p 0.672904mV 990102.144p 0.672904mV 990115.685p 0.686234mV 990134.276p 0.725543mV 991016.369p 0.58125mV 992053.487p 0.68623mV 992077.126p 0.736357mV 993027.629p 0.475374mV 993043.113p 0.444355mV 993053.324p 0.418695mV 993056.471p 0.401648mV 993057.886p 0.401648mV 994056.972p 0.335031mV 995029.183p 0.528272mV 995058.268p 0.350258mV 996007.06p 0.598422mV 996018.075p 0.618448mV 996021.251p 0.625816mV 996047.063p 0.650947mV 996049.149p 0.650947mV 996081.092p 0.655156mV 996095.212p 0.738395mV 997020.477p 0.574466mV 997021.648p 0.574466mV 997033.211p 0.581504mV 997066.838p 0.494272mV 997081.206p 0.395127mV 998002.499p 0.52461mV 998015.241p 0.527804mV 998068.603p 0.708829mV 998076.926p 0.754884mV 999001.686p 0.502096mV 999061.006p 0.416985mV)
.ENDS conductors__anyBias-Lk_0_703

.SUBCKT conductors__anyBias-Lk_0_704 bottom out
VrampSppl@0 bottom out pwl(0 0 1001.357p 0.546987mV 1003.807p 0.546987mV 1033.68p 0.442384mV 1057.776p 0.403003mV 2026.674p 0.574766mV 2103.161p 0.502997mV 2117.296p 0.423717mV 3014.209p 0.54801mV 3022.9p 0.598174mV 3028.376p 0.623402mV 3040.213p 0.595927mV 4002.784p 0.547468mV 4012.055p 0.550015mV 4035.68p 0.636103mV 4046.911p 0.693985mV 5053.928p 0.58983mV 5121.883p 0.711606mV 6009.897p 0.520153mV 6011.833p 0.494569mV 6037.964p 0.574237mV 6042.09p 0.600404mV 6070.71p 0.712492mV 7011.005p 0.605675mV 7017.232p 0.580941mV 7027.676p 0.584975mV 7033.505p 0.61368mV 7049.208p 0.544322mV 7052.476p 0.573896mV 7052.928p 0.573896mV 7059.424p 0.551194mV 7105.76p 0.637934mV 7117.36p 0.645544mV 8044.351p 0.543479mV 8047.479p 0.51539mV 8053.171p 0.53982mV 8056.57p 0.564015mV 8070.528p 0.584314mV 8083.563p 0.633635mV 8084.332p 0.633635mV 8118.998p 0.664908mV 9005.414p 0.524971mV 10008.846p 0.577029mV 10017.442p 0.627654mV 10018.242p 0.627654mV 10024.941p 0.653395mV 10032.688p 0.706508mV 10034.526p 0.706508mV 10037.457p 0.681546mV 10043.297p 0.710109mV 10051.973p 0.717224mV 10052.398p 0.717224mV 10054.04p 0.717224mV 11015.92p 0.524636mV 11029.904p 0.526031mV 11035.681p 0.473789mV 12047.943p 0.586345mV 12062.291p 0.571388mV 12075.402p 0.609473mV 12093.636p 0.650412mV 13039.024p 0.579374mV 13057.94p 0.636033mV 13062.288p 0.664057mV 13099.399p 0.611296mV 13108.489p 0.672643mV 14057.256p 0.64332mV 14075.153p 0.603742mV 15003.841p 0.547695mV 15018.256p 0.575726mV 15068.18p 0.645483mV 15083.34p 0.682672mV 16032.353p 0.593741mV 16036.351p 0.618532mV 16045.204p 0.669144mV 16051.409p 0.695275mV 16054.411p 0.695275mV 16064.298p 0.644614mV 16069.417p 0.62056mV 17004.853p 0.548995mV 17049.718p 0.507757mV 18015.66p 0.630509mV 18026.594p 0.631976mV 18055.949p 0.541844mV 18069.821p 0.600948mV 18074.743p 0.578378mV 18095.434p 0.626222mV 18098.778p 0.626222mV 19004.144p 0.549136mV 19025.369p 0.624271mV 19027.509p 0.624271mV 19036.73p 0.57146mV 19043.36p 0.598267mV 19051.564p 0.599786mV 19076.379p 0.635791mV 20025.27p 0.581426mV 20029.434p 0.581426mV 20038.146p 0.637979mV 21004.905p 0.549697mV 21031.907p 0.547791mV 21034.558p 0.547791mV 21055.108p 0.468857mV 21082.246p 0.382238mV 22040.469p 0.550673mV 22043.173p 0.550673mV 22046.205p 0.57801mV 22063.074p 0.660693mV 22072.375p 0.613032mV 22127.179p 0.413117mV 22140.614p 0.385692mV 23046.135p 0.620615mV 23062.198p 0.646107mV 23071.34p 0.595021mV 23095.069p 0.738258mV 24009.38p 0.518984mV 25010.159p 0.551293mV 25015.533p 0.576892mV 25065.559p 0.569823mV 25095.767p 0.56142mV 25115.141p 0.610205mV 25119.908p 0.610205mV 25138.179p 0.718476mV 25143.871p 0.694751mV 26018.557p 0.467462mV 26024.846p 0.49361mV 26031.56p 0.54448mV 26038.005p 0.516905mV 26081.853p 0.528843mV 26103.278p 0.468642mV 26119.938p 0.432494mV 27008.06p 0.526071mV 27016.641p 0.475011mV 27022.32p 0.501761mV 27022.633p 0.501761mV 27037.914p 0.4745mV 27045.765p 0.419774mV 27048.114p 0.419774mV 27065.969p 0.460231mV 28009.804p 0.523837mV 28024.494p 0.552659mV 28029.225p 0.579401mV 28041.218p 0.502047mV 29037.282p 0.417401mV 29052.261p 0.38572mV 30015.036p 0.528572mV 30058.187p 0.525303mV 30094.296p 0.585407mV 30102.965p 0.63167mV 30103.588p 0.63167mV 30111.938p 0.627035mV 30117.433p 0.651958mV 30148.117p 0.656455mV 30159.327p 0.663377mV 30161.043p 0.642027mV 31064.957p 0.503091mV 31084.216p 0.501757mV 31089.256p 0.52649mV 31102.229p 0.441495mV 31113.594p 0.487463mV 31129.812p 0.447897mV 32053.048p 0.588848mV 32065.331p 0.666617mV 32071.652p 0.640785mV 32076.459p 0.615711mV 32078.883p 0.615711mV 32079.463p 0.615711mV 32081.237p 0.643802mV 32092.176p 0.648773mV 32092.241p 0.648773mV 32105.136p 0.738575mV 33005.182p 0.528572mV 33016.401p 0.52947mV 33049.011p 0.527688mV 33056.041p 0.526461mV 33092.762p 0.65359mV 33093.114p 0.65359mV 33098.746p 0.681216mV 33107.573p 0.686008mV 33114.9p 0.715835mV 34022.666p 0.543922mV 34035.994p 0.565976mV 34037.451p 0.565976mV 34042.225p 0.538582mV 34051.972p 0.589209mV 34058.18p 0.561928mV 34065.433p 0.560586mV 34110.458p 0.466771mV 34118.874p 0.48919mV 34148.243p 0.563618mV 34156.999p 0.604417mV 34227.935p 0.622539mV 34242.981p 0.600618mV 34260.051p 0.662492mV 34271.994p 0.669853mV 35027.603p 0.520071mV 35074.82p 0.522191mV 35081.94p 0.512233mV 35094.088p 0.501802mV 36011.784p 0.596865mV 36037.184p 0.622722mV 36053.155p 0.6015mV 36067.079p 0.635097mV 37016.167p 0.577043mV 37033.151p 0.601967mV 37076.303p 0.69485mV 38047.848p 0.577605mV 38064.102p 0.607639mV 38075.005p 0.640285mV 39031.725p 0.555129mV 39031.821p 0.555129mV 39034.508p 0.555129mV 39044.902p 0.556839mV 39065.492p 0.534756mV 39076.762p 0.482032mV 39096.537p 0.531457mV 39099.869p 0.531457mV 39126.861p 0.517825mV 39149.778p 0.501866mV 39150.487p 0.523107mV 39155.071p 0.543992mV 40001.855p 0.546636mV 40010.453p 0.548424mV 40013.223p 0.548424mV 40018.456p 0.523137mV 40033.54p 0.499211mV 40052.271p 0.552114mV 40081.721p 0.500527mV 40137.291p 0.562132mV 40140.126p 0.585754mV 40182.43p 0.624694mV 40192.137p 0.571629mV 40213.281p 0.573504mV 40218.437p 0.600736mV 40220.115p 0.575468mV 40225.959p 0.550535mV 40234.424p 0.525772mV 40239.301p 0.553606mV 40241.378p 0.581297mV 40245.124p 0.609008mV 40247.935p 0.609008mV 41006.777p 0.580514mV 41023.288p 0.556245mV 41102.626p 0.628548mV 42007.856p 0.581396mV 42047.824p 0.656168mV 42048.28p 0.656168mV 42053.892p 0.635272mV 42054.697p 0.635272mV 43003.362p 0.551271mV 43024.727p 0.547165mV 43027.341p 0.572189mV 43040.809p 0.489582mV 43052.68p 0.486417mV 43062.594p 0.534503mV 43063.436p 0.534503mV 43097.874p 0.536981mV 43158.291p 0.592328mV 43169.809p 0.638784mV 43170.007p 0.662616mV 43199.107p 0.633746mV 43211.195p 0.71905mV 44016.337p 0.629657mV 44026.593p 0.631127mV 44029.464p 0.631127mV 44045.531p 0.640395mV 45019.266p 0.471142mV 45030.299p 0.543871mV 45060.082p 0.419311mV 46033.335p 0.549777mV 46034.917p 0.549777mV 46040.846p 0.603488mV 46058.306p 0.580435mV 46066.543p 0.636914mV 46072.066p 0.613112mV 47014.887p 0.546905mV 47029.21p 0.519127mV 47032.833p 0.492156mV 47083.776p 0.58639mV 47089.517p 0.612386mV 47090.412p 0.638614mV 47093.389p 0.638614mV 47094.856p 0.638614mV 47108.98p 0.615mV 47138.49p 0.632029mV 48016.558p 0.464255mV 48017.801p 0.464255mV 49057.74p 0.50728mV 49061.493p 0.530758mV 50042.417p 0.49395mV 50045.738p 0.519735mV 50049.557p 0.519735mV 50051.866p 0.492505mV 50081.142p 0.53594mV 50093.67p 0.584569mV 50110.93p 0.631343mV 50112.311p 0.631343mV 50143.327p 0.638271mV 50156.229p 0.623961mV 50156.884p 0.623961mV 50185.693p 0.553081mV 50190.261p 0.584363mV 50194.946p 0.584363mV 50201.41p 0.595592mV 51006.115p 0.519196mV 51065.941p 0.608049mV 51077.848p 0.607016mV 51089.024p 0.555094mV 51115.114p 0.614795mV 51133.17p 0.595146mV 52013.694p 0.549671mV 52024.012p 0.496926mV 52037.555p 0.52183mV 52051.188p 0.492674mV 52065.832p 0.460823mV 52066.129p 0.460823mV 53014.646p 0.603336mV 53016.744p 0.578518mV 53067.218p 0.552734mV 53074.307p 0.582567mV 54006.263p 0.527272mV 54010.924p 0.55332mV 54016.49p 0.579222mV 54067.896p 0.696058mV 54068.542p 0.696058mV 54071.682p 0.725808mV 55004.023p 0.545792mV 55025.951p 0.46244mV 55030.703p 0.486388mV 56034.78p 0.500158mV 56049.914p 0.524652mV 56052.088p 0.497195mV 56055.382p 0.522207mV 56056.537p 0.522207mV 56056.598p 0.522207mV 56081.785p 0.538108mV 56084.552p 0.538108mV 56089.334p 0.509572mV 56097.21p 0.504608mV 57031.129p 0.611749mV 57068.492p 0.609611mV 58037.523p 0.476509mV 58057.84p 0.578375mV 58058.781p 0.578375mV 58112.181p 0.481034mV 59059.338p 0.464649mV 59075.996p 0.451489mV 59076.936p 0.451489mV 59083.118p 0.421236mV 60033.466p 0.5043mV 60039.743p 0.53026mV 60070.233p 0.551299mV 60074.607p 0.551299mV 60112.258p 0.71435mV 60118.756p 0.743953mV 61011.898p 0.552294mV 61035.973p 0.583816mV 61109.387p 0.502571mV 61156.462p 0.54592mV 61159.852p 0.54592mV 61180.254p 0.563448mV 61209.349p 0.529607mV 61220.02p 0.445976mV 61221.412p 0.445976mV 61232.095p 0.440798mV 61237.799p 0.463476mV 62028.202p 0.5717mV 62054.658p 0.600464mV 62090.623p 0.566358mV 62126.681p 0.567238mV 62143.75p 0.606393mV 63031.749p 0.547865mV 63036.952p 0.57338mV 63042.965p 0.546224mV 63049.575p 0.571877mV 63128.918p 0.455278mV 63134.963p 0.479286mV 64008.948p 0.523086mV 64016.084p 0.52364mV 66002.813p 0.55085mV 66039.614p 0.471393mV 66057.104p 0.514288mV 66061.624p 0.536974mV 66071.356p 0.581743mV 67007.742p 0.525563mV 67008.567p 0.525563mV 67037.83p 0.462367mV 68000.065p 0.553516mV 68001.766p 0.553516mV 68002.988p 0.553516mV 68044.862p 0.492593mV 68068.294p 0.497703mV 69009.777p 0.580214mV 69036.891p 0.536792mV 69039.58p 0.536792mV 69084.202p 0.469861mV 69096.014p 0.441231mV 69112.828p 0.511266mV 69115.605p 0.481387mV 69115.985p 0.481387mV 69134.602p 0.494094mV 70044.898p 0.610086mV 70060.128p 0.673728mV 70060.19p 0.673728mV 70061.559p 0.673728mV 71007.717p 0.579696mV 71017.333p 0.527413mV 71026.879p 0.475218mV 71031.111p 0.501425mV 71040.414p 0.447248mV 71044.738p 0.447248mV 72000.556p 0.545793mV 72017.61p 0.569793mV 72032.469p 0.594132mV 72034.073p 0.594132mV 72046.796p 0.566848mV 72046.918p 0.566848mV 72050.098p 0.540297mV 72094.307p 0.652104mV 72102.168p 0.659448mV 72104.822p 0.659448mV 72105.356p 0.689915mV 73013.833p 0.552202mV 73025.353p 0.523496mV 73060.297p 0.540844mV 73064.558p 0.540844mV 73079.947p 0.559329mV 73131.339p 0.66066mV 73170.184p 0.554748mV 73176.494p 0.581578mV 73184.101p 0.555763mV 73202.876p 0.612191mV 75053.123p 0.541388mV 75091.777p 0.532276mV 75095.914p 0.504146mV 75103.021p 0.528452mV 75111.258p 0.576292mV 75115.571p 0.547685mV 75123.313p 0.571727mV 75134.111p 0.514911mV 75177.457p 0.631685mV 75187.947p 0.68686mV 75192.402p 0.662816mV 76052.704p 0.453609mV 76083.788p 0.549955mV 76092.418p 0.598286mV 76093.513p 0.598286mV 76111.384p 0.53997mV 76172.201p 0.541558mV 76186.27p 0.568598mV 76187.426p 0.568598mV 76192.786p 0.542278mV 76233.033p 0.596714mV 76258.394p 0.687325mV 77016.411p 0.580676mV 77033.884p 0.504221mV 77044.74p 0.505538mV 77087.284p 0.51391mV 78004.035p 0.550454mV 78030.08p 0.61314mV 78050.71p 0.677723mV 78054.352p 0.677723mV 79006.408p 0.578088mV 79006.547p 0.578088mV 79024.086p 0.556261mV 79048.788p 0.589854mV 79068.907p 0.597895mV 79084.638p 0.684888mV 79088.286p 0.7148mV 80025.031p 0.618887mV 80046.059p 0.618753mV 80050.036p 0.646191mV 80053.869p 0.646191mV 80074.558p 0.656953mV 80075.937p 0.687542mV 80076.885p 0.687542mV 81136.929p 0.550865mV 81143.4p 0.575904mV 81149.915p 0.548326mV 81156.514p 0.546109mV 81195.047p 0.594005mV 81208.466p 0.64765mV 81221.711p 0.573673mV 81257.127p 0.619065mV 81277.439p 0.582646mV 81284.344p 0.613395mV 82004.187p 0.552736mV 82062.653p 0.564085mV 82073.996p 0.567602mV 82079.288p 0.595625mV 82083.033p 0.571196mV 82083.511p 0.571196mV 82090.668p 0.575611mV 82098.688p 0.604408mV 82107.009p 0.557863mV 82109.043p 0.557863mV 82140.129p 0.447848mV 82210.086p 0.444514mV 82240.469p 0.471679mV 82241.764p 0.471679mV 83016.041p 0.46809mV 83022.812p 0.494374mV 83038.807p 0.465085mV 83062.808p 0.476535mV 83062.884p 0.476535mV 84015.49p 0.522272mV 84047.181p 0.412747mV 85030.332p 0.546874mV 85079.222p 0.515667mV 85086.876p 0.511257mV 86027.152p 0.575554mV 86030.345p 0.549812mV 86058.73p 0.634276mV 86065.434p 0.639743mV 86074.402p 0.617333mV 86080.942p 0.626286mV 86087.564p 0.657354mV 87065.225p 0.698501mV 88040.552p 0.58371mV 88097.17p 0.543426mV 88103.044p 0.515385mV 88130.29p 0.607403mV 88143.661p 0.656035mV 88165.689p 0.789463mV 89021.674p 0.440712mV 89023.903p 0.440712mV 90000.304p 0.546856mV 90061.88p 0.560036mV 90082.568p 0.461783mV 90131.42p 0.452465mV 91001.373p 0.549201mV 91013.374p 0.49699mV 91028.996p 0.522682mV 91033.472p 0.495577mV 91060.929p 0.589595mV 91084.44p 0.634928mV 92005.287p 0.576953mV 92015.235p 0.524045mV 92021.566p 0.497678mV 92045.649p 0.412861mV 92055.689p 0.353527mV 93012.727p 0.494329mV 93015.089p 0.467812mV 93023.59p 0.493622mV 94019.916p 0.526336mV 94063.6p 0.479961mV 94064.549p 0.479961mV 94068.734p 0.502011mV 94096.413p 0.576181mV 94106.411p 0.565958mV 94109.476p 0.565958mV 94117.728p 0.555921mV 94133.026p 0.566833mV 94139.369p 0.536048mV 94152.837p 0.599246mV 94175.456p 0.447279mV 94180.326p 0.416425mV 95013.897p 0.604375mV 95069.716p 0.652772mV 96010.487p 0.605307mV 96016.022p 0.63301mV 96020.446p 0.661036mV 96025.715p 0.637045mV 96029.775p 0.637045mV 96034.0p 0.613823mV 96036.963p 0.591217mV 96045.928p 0.599246mV 96060.87p 0.586844mV 96076.539p 0.575857mV 97000.233p 0.554285mV 97073.077p 0.545597mV 97119.971p 0.554849mV 97123.138p 0.527003mV 97126.697p 0.551782mV 97129.166p 0.551782mV 97129.259p 0.551782mV 97140.104p 0.467793mV 97163.014p 0.404176mV 98001.354p 0.546625mV 98018.999p 0.571716mV 98033.073p 0.651246mV 98045.518p 0.629748mV 98045.733p 0.629748mV 99012.689p 0.603482mV 99049.189p 0.688349mV 100015.201p 0.629919mV 100017.602p 0.629919mV 100028.296p 0.630207mV 100058.161p 0.64228mV 100068.976p 0.598231mV 101002.399p 0.547021mV 101017.086p 0.521287mV 101020.378p 0.547686mV 101084.64p 0.525487mV 101096.477p 0.537191mV 101129.598p 0.507202mV 102017.333p 0.530291mV 102063.388p 0.451665mV 103006.456p 0.576127mV 103008.329p 0.576127mV 104005.47p 0.525367mV 104016.046p 0.575576mV 104019.771p 0.575576mV 104068.351p 0.52062mV 104083.602p 0.546518mV 104095.049p 0.571728mV 104119.845p 0.57061mV 104125.247p 0.517177mV 104128.05p 0.517177mV 104195.232p 0.572446mV 104220.35p 0.555167mV 104251.254p 0.617997mV 104261.222p 0.623965mV 104292.389p 0.549365mV 104293.327p 0.549365mV 104343.111p 0.552134mV 104357.427p 0.54303mV 105011.412p 0.548986mV 105034.047p 0.546847mV 105036.028p 0.572528mV 105042.3p 0.598189mV 105050.54p 0.59743mV 105073.868p 0.547202mV 105078.609p 0.522004mV 105083.229p 0.549426mV 105085.743p 0.524027mV 106018.194p 0.521202mV 106045.163p 0.465947mV 106051.068p 0.491179mV 107030.706p 0.497187mV 107041.521p 0.547173mV 107049.406p 0.519225mV 107051.911p 0.54384mV 107073.137p 0.535759mV 107115.198p 0.589597mV 107122.167p 0.560309mV 107169.137p 0.619573mV 107188.857p 0.673273mV 107208.909p 0.579952mV 107223.303p 0.618776mV 107229.329p 0.649499mV 108006.156p 0.580601mV 108018.128p 0.58211mV 108038.246p 0.692739mV 108040.869p 0.66923mV 108047.838p 0.646724mV 109014.099p 0.495352mV 110008.495p 0.523333mV 110016.513p 0.523476mV 110035.759p 0.520378mV 110055.91p 0.565301mV 110077.012p 0.503957mV 110080.152p 0.527645mV 110083.793p 0.527645mV 111001.335p 0.554343mV 111057.928p 0.575291mV 111069.959p 0.521479mV 111073.915p 0.49464mV 111080.645p 0.440278mV 111084.968p 0.440278mV 112010.845p 0.546686mV 112022.044p 0.49451mV 112037.532p 0.467135mV 112054.223p 0.435678mV 113016.704p 0.58214mV 113046.377p 0.483186mV 113080.551p 0.402007mV 114008.897p 0.574491mV 114035.314p 0.516155mV 114035.886p 0.516155mV 114045.805p 0.51278mV 114061.16p 0.584408mV 114062.203p 0.584408mV 114068.539p 0.608213mV 114090.778p 0.573785mV 114142.059p 0.62656mV 114158.798p 0.714467mV 114161.654p 0.693069mV 115047.777p 0.538956mV 115071.786p 0.679799mV 116027.25p 0.575935mV 116036.852p 0.628213mV 116049.718p 0.576447mV 116065.348p 0.634905mV 116067.369p 0.634905mV 116068.935p 0.634905mV 116072.376p 0.611424mV 116095.169p 0.552251mV 116100.49p 0.530701mV 116110.543p 0.539432mV 116123.594p 0.600104mV 117043.057p 0.653349mV 118053.553p 0.712351mV 119004.709p 0.54718mV 119036.029p 0.563937mV 119046.6p 0.560354mV 119071.998p 0.471593mV 119091.858p 0.457711mV 120005.521p 0.573899mV 120017.449p 0.57599mV 120022.059p 0.551128mV 120030.405p 0.606931mV 120032.934p 0.606931mV 120056.988p 0.699752mV 120057.958p 0.699752mV 121009.007p 0.52433mV 121016.309p 0.471107mV 121065.17p 0.495329mV 122003.727p 0.547327mV 122004.737p 0.547327mV 122052.79p 0.490619mV 122072.137p 0.527809mV 122083.339p 0.466534mV 123005.848p 0.521175mV 123015.628p 0.520053mV 123026.216p 0.518515mV 123044.01p 0.435197mV 124013.27p 0.603891mV 124064.802p 0.624743mV 125000.085p 0.547399mV 125016.656p 0.469893mV 125043.9p 0.491021mV 125045.008p 0.515087mV 125049.674p 0.515087mV 126007.464p 0.52262mV 126016.895p 0.523089mV 126019.093p 0.523089mV 126043.022p 0.549122mV 126076.196p 0.465868mV 126077.368p 0.465868mV 126096.832p 0.453329mV 126097.198p 0.453329mV 126107.416p 0.443939mV 127028.897p 0.629223mV 127062.492p 0.67895mV 128048.784p 0.691866mV 128050.29p 0.669721mV 129036.109p 0.468267mV 129044.457p 0.440638mV 130008.95p 0.522291mV 130039.121p 0.529509mV 130098.817p 0.537396mV 130103.443p 0.509993mV 130117.984p 0.532227mV 130141.933p 0.656979mV 130143.024p 0.656979mV 130154.009p 0.656777mV 130158.175p 0.683843mV 130160.63p 0.711545mV 130165.429p 0.68752mV 130177.482p 0.694932mV 131034.482p 0.604597mV 131037.266p 0.578977mV 131125.551p 0.465641mV 132007.916p 0.579178mV 132008.375p 0.579178mV 132027.407p 0.523932mV 132080.609p 0.52776mV 132116.856p 0.584606mV 132117.773p 0.584606mV 132148.781p 0.572546mV 132178.976p 0.617662mV 132181.308p 0.590957mV 132208.472p 0.565851mV 132238.773p 0.675835mV 132243.643p 0.704531mV 132247.168p 0.681628mV 132251.197p 0.711832mV 134006.664p 0.527054mV 134006.779p 0.527054mV 134012.096p 0.501974mV 134028.364p 0.47784mV 134076.497p 0.507004mV 135000.022p 0.551394mV 135000.209p 0.551394mV 135008.739p 0.526291mV 135019.643p 0.528575mV 135033.732p 0.505299mV 135034.7p 0.505299mV 135035.351p 0.479846mV 135073.256p 0.395444mV 136007.959p 0.520145mV 136042.608p 0.53494mV 136075.073p 0.649626mV 136084.064p 0.675279mV 136091.547p 0.675945mV 136094.909p 0.675945mV 136095.104p 0.650985mV 136097.955p 0.650985mV 136100.196p 0.626869mV 136123.946p 0.693704mV 137038.105p 0.569943mV 137093.179p 0.606022mV 138008.79p 0.573076mV 138011.796p 0.547097mV 138028.269p 0.522059mV 138055.561p 0.519841mV 138099.618p 0.606992mV 138124.957p 0.572129mV 138125.976p 0.544999mV 138126.766p 0.544999mV 138144.907p 0.516747mV 138160.204p 0.512346mV 138167.721p 0.536471mV 138187.446p 0.420974mV 138192.855p 0.443297mV 139007.204p 0.523286mV 139067.049p 0.562505mV 139100.903p 0.474894mV 139101.212p 0.474894mV 139115.277p 0.439466mV 139117.366p 0.439466mV 139120.548p 0.461524mV 140036.179p 0.474274mV 141027.834p 0.582549mV 141048.301p 0.537164mV 141050.241p 0.565531mV 141075.671p 0.497348mV 141079.296p 0.497348mV 141090.258p 0.475861mV 141098.871p 0.503049mV 141100.017p 0.529782mV 141112.042p 0.582536mV 141116.82p 0.556206mV 141156.56p 0.55946mV 141170.019p 0.536877mV 141198.3p 0.517555mV 141202.464p 0.492866mV 141233.366p 0.439997mV 142019.076p 0.577387mV 142019.728p 0.577387mV 142028.803p 0.579413mV 142044.156p 0.609817mV 143009.691p 0.576521mV 143036.612p 0.627894mV 144005.576p 0.521159mV 144041.958p 0.550498mV 144045.886p 0.578222mV 144046.255p 0.578222mV 144053.215p 0.553341mV 144063.478p 0.556563mV 144074.612p 0.559577mV 144083.368p 0.615069mV 144085.389p 0.590487mV 144111.424p 0.62862mV 144132.838p 0.643372mV 145002.331p 0.546057mV 145003.919p 0.546057mV 145009.978p 0.519219mV 145024.066p 0.490568mV 145033.305p 0.435032mV 145033.791p 0.435032mV 145048.677p 0.452151mV 145053.882p 0.473553mV 146005.811p 0.524293mV 146011.949p 0.549321mV 146036.713p 0.569589mV 146058.608p 0.567075mV 146101.095p 0.48237mV 146112.415p 0.476929mV 146133.179p 0.407931mV 147000.162p 0.553823mV 147030.208p 0.599245mV 147032.459p 0.599245mV 147042.889p 0.597173mV 147048.508p 0.622754mV 147080.341p 0.651037mV 148034.604p 0.612994mV 148043.851p 0.617595mV 148058.233p 0.705693mV 149016.644p 0.523086mV 149038.04p 0.474083mV 149107.305p 0.537943mV 150051.962p 0.493555mV 150066.398p 0.462184mV 150070.948p 0.485867mV 150078.527p 0.508937mV 150085.092p 0.501662mV 151063.006p 0.419036mV 152016.549p 0.528885mV 152021.67p 0.504073mV 153005.788p 0.523422mV 153053.481p 0.474636mV 154003.193p 0.547704mV 154004.009p 0.547704mV 154024.798p 0.552734mV 154078.812p 0.593955mV 154080.389p 0.569491mV 154095.545p 0.602231mV 154103.271p 0.630803mV 154118.987p 0.666563mV 155008.5p 0.57314mV 155032.252p 0.551963mV 155055.483p 0.586409mV 155078.658p 0.702967mV 156031.151p 0.506998mV 156033.011p 0.506998mV 156066.262p 0.479113mV 156100.079p 0.427497mV 157024.574p 0.606409mV 157044.045p 0.719419mV 158007.473p 0.57668mV 158023.879p 0.660351mV 158045.94p 0.652582mV 159017.687p 0.469017mV 159024.176p 0.493767mV 159024.624p 0.493767mV 159032.04p 0.489323mV 159047.451p 0.401712mV 160003.228p 0.548631mV 160019.406p 0.574868mV 160020.783p 0.601596mV 160028.501p 0.575806mV 160029.978p 0.575806mV 160046.451p 0.580634mV 160047.244p 0.580634mV 160048.75p 0.580634mV 160055.631p 0.584595mV 160065.194p 0.589072mV 160087.449p 0.601158mV 161051.156p 0.601873mV 161056.076p 0.575713mV 161073.243p 0.551225mV 161087.772p 0.579937mV 161134.549p 0.455025mV 161148.063p 0.476652mV 161171.822p 0.592646mV 161178.544p 0.563317mV 161186.686p 0.609946mV 161190.948p 0.633564mV 161197.484p 0.605099mV 161214.702p 0.680131mV 162001.163p 0.547955mV 163015.476p 0.575269mV 163032.78p 0.551126mV 163041.915p 0.4997mV 163046.453p 0.526507mV 163075.647p 0.472867mV 163094.72p 0.389669mV 163104.906p 0.382914mV 164000.155p 0.548708mV 164008.313p 0.521334mV 164020.036p 0.491105mV 164029.783p 0.515246mV 164057.431p 0.442608mV 165029.561p 0.465568mV 166000.818p 0.546808mV 166007.777p 0.574338mV 167027.905p 0.687516mV 168018.923p 0.470324mV 169029.032p 0.474256mV 169063.645p 0.545375mV 169068.899p 0.569713mV 169093.285p 0.48053mV 169127.63p 0.530884mV 169140.463p 0.489923mV 170016.716p 0.523176mV 170027.936p 0.525104mV 170064.543p 0.444395mV 172001.545p 0.547534mV 172039.358p 0.516258mV 172059.945p 0.563092mV 172060.914p 0.5349mV 172065.508p 0.506785mV 172077.188p 0.450135mV 172086.885p 0.444301mV 172108.401p 0.426341mV 173020.084p 0.596718mV 173025.36p 0.569891mV 173050.726p 0.489469mV 173052.333p 0.489469mV 173059.817p 0.461919mV 174014.646p 0.598652mV 174043.54p 0.540634mV 174071.709p 0.483mV 174073.124p 0.483mV 174087.903p 0.503414mV 174178.959p 0.535311mV 174183.678p 0.505004mV 174200.535p 0.536868mV 175010.184p 0.497368mV 176045.381p 0.639134mV 176057.559p 0.592685mV 176062.399p 0.622422mV 176069.312p 0.652379mV 177041.682p 0.478331mV 177046.227p 0.448875mV 178005.233p 0.576431mV 178007.725p 0.576431mV 178009.288p 0.576431mV 178030.513p 0.491608mV 179003.529p 0.551528mV 179022.091p 0.657725mV 179039.614p 0.688983mV 179047.603p 0.747915mV 180013.459p 0.554921mV 180018.96p 0.581954mV 180040.255p 0.560016mV 180090.656p 0.581969mV 180111.11p 0.649209mV 180111.152p 0.649209mV 181009.907p 0.521923mV 181013.271p 0.548914mV 181033.24p 0.497798mV 181035.14p 0.471596mV 181049.066p 0.470729mV 181051.543p 0.49604mV 181053.441p 0.49604mV 181066.533p 0.516949mV 181069.036p 0.516949mV 181082.466p 0.589023mV 181134.008p 0.632718mV 182051.454p 0.620007mV 183066.446p 0.584544mV 183077.164p 0.638911mV 183099.078p 0.594447mV 183111.531p 0.52457mV 183112.434p 0.52457mV 183152.612p 0.48599mV 183154.767p 0.48599mV 183155.376p 0.458896mV 183165.578p 0.456025mV 184009.242p 0.52587mV 184066.06p 0.569413mV 184067.001p 0.569413mV 184073.398p 0.595995mV 184083.805p 0.544341mV 184095.242p 0.572752mV 184141.097p 0.499436mV 185005.619p 0.519506mV 185015.253p 0.519334mV 185028.086p 0.570727mV 185069.585p 0.507299mV 186009.184p 0.576109mV 186030.871p 0.503255mV 186047.704p 0.425542mV 186056.321p 0.423574mV 186056.704p 0.423574mV 187004.965p 0.553479mV 187021.193p 0.603228mV 187021.751p 0.603228mV 187025.394p 0.576686mV 187032.917p 0.60316mV 187043.204p 0.656771mV 187065.95p 0.748167mV 188038.964p 0.457383mV 189009.404p 0.57757mV 189038.866p 0.464217mV 189040.722p 0.435808mV 190005.789p 0.525591mV 190032.356p 0.557098mV 190048.773p 0.53425mV 190050.226p 0.508742mV 190065.823p 0.536629mV 190068.117p 0.536629mV 190096.98p 0.591798mV 190107.766p 0.593023mV 190110.064p 0.620198mV 190112.339p 0.620198mV 190136.725p 0.656229mV 190151.264p 0.64324mV 191006.572p 0.52067mV 191028.104p 0.461396mV 192015.481p 0.518169mV 192030.652p 0.539521mV 192057.292p 0.555401mV 192058.225p 0.555401mV 192073.482p 0.520893mV 192086.42p 0.537105mV 192090.557p 0.507671mV 192094.326p 0.507671mV 192102.076p 0.500689mV 192122.428p 0.484042mV 193033.149p 0.438996mV 193054.706p 0.426658mV 193059.157p 0.396065mV 194025.573p 0.634551mV 194026.75p 0.634551mV 194057.204p 0.60359mV 194064.187p 0.634725mV 195003.616p 0.551469mV 195045.56p 0.628962mV 195063.874p 0.556248mV 195066.016p 0.58507mV 195094.854p 0.626527mV 196066.066p 0.498364mV 197000.267p 0.548668mV 197018.686p 0.519735mV 197030.232p 0.541614mV 197034.482p 0.541614mV 197047.17p 0.458076mV 197051.53p 0.482221mV 197053.371p 0.482221mV 197075.388p 0.544436mV 197086.483p 0.537658mV 198098.639p 0.59853mV 199006.938p 0.522311mV 199037.717p 0.568712mV 199064.974p 0.536084mV 199114.013p 0.456467mV 200012.01p 0.54561mV 200026.852p 0.518386mV 200057.885p 0.457969mV 200061.22p 0.481628mV 200083.51p 0.467223mV 200085.808p 0.488901mV 201023.846p 0.609852mV 201031.65p 0.665634mV 201040.797p 0.618609mV 201058.874p 0.656565mV 201058.883p 0.656565mV 202026.079p 0.522045mV 202048.605p 0.467115mV 202049.331p 0.467115mV 202075.671p 0.450106mV 203015.21p 0.53072mV 203031.388p 0.614179mV 203058.132p 0.651845mV 203061.149p 0.681201mV 204019.948p 0.524226mV 204025.292p 0.469328mV 204052.08p 0.428206mV 205033.952p 0.593699mV 205062.141p 0.647744mV 205064.349p 0.647744mV 205065.997p 0.67601mV 205086.802p 0.690863mV 206038.755p 0.523422mV 206075.427p 0.518008mV 206085.25p 0.460928mV 206088.16p 0.460928mV 206090.827p 0.484356mV 207017.425p 0.582951mV 207039.128p 0.588045mV 207066.879p 0.602342mV 207099.402p 0.628882mV 208006.428p 0.520247mV 208012.164p 0.545242mV 208047.892p 0.561576mV 208065.87p 0.609611mV 208066.033p 0.609611mV 208068.157p 0.609611mV 208078.083p 0.662325mV 209018.372p 0.57474mV 209028.172p 0.576551mV 209030.18p 0.551208mV 209030.583p 0.551208mV 209047.495p 0.528195mV 209091.029p 0.451888mV 210007.797p 0.529226mV 210021.999p 0.506703mV 210051.006p 0.511526mV 210058.258p 0.537949mV 210089.922p 0.587471mV 210093.904p 0.560327mV 210094.876p 0.560327mV 210108.12p 0.532607mV 210141.85p 0.55271mV 210148.892p 0.52454mV 210180.432p 0.532589mV 210188.56p 0.555613mV 210226.03p 0.472753mV 211021.722p 0.544484mV 211047.35p 0.514379mV 211059.885p 0.511981mV 211068.352p 0.561575mV 211124.001p 0.51728mV 211132.421p 0.460597mV 211135.237p 0.431821mV 211138.669p 0.431821mV 212013.118p 0.606256mV 212017.761p 0.633216mV 212064.293p 0.580044mV 212075.956p 0.620341mV 213008.899p 0.526052mV 213030.129p 0.492075mV 213036.605p 0.516204mV 213057.711p 0.504583mV 213070.136p 0.467079mV 214007.303p 0.519972mV 214023.037p 0.43761mV 214036.0p 0.350914mV 215023.752p 0.49822mV 215033.65p 0.497664mV 215053.129p 0.544858mV 215075.408p 0.507018mV 215122.953p 0.552634mV 215144.323p 0.536413mV 215163.76p 0.466385mV 215166.055p 0.435248mV 216023.289p 0.595782mV 216032.287p 0.594347mV 216043.939p 0.59371mV 216082.52p 0.598316mV 216085.392p 0.626742mV 217012.657p 0.548784mV 217014.056p 0.548784mV 218026.681p 0.62041mV 218053.336p 0.649935mV 218069.133p 0.684646mV 219001.917p 0.547297mV 219013.86p 0.54978mV 219020.469p 0.499254mV 219044.366p 0.447609mV 219044.88p 0.447609mV 219049.899p 0.472568mV 219053.529p 0.444308mV 220054.447p 0.534364mV 220073.505p 0.57754mV 220092.514p 0.620496mV 220116.377p 0.642984mV 220122.627p 0.618188mV 220140.119p 0.734435mV 220143.49p 0.734435mV 221007.108p 0.523474mV 221055.099p 0.524781mV 221055.84p 0.524781mV 221061.219p 0.550073mV 221061.748p 0.550073mV 221077.346p 0.572979mV 221083.024p 0.5986mV 221106.224p 0.518132mV 221124.777p 0.542529mV 221128.908p 0.567684mV 221131.872p 0.592789mV 221141.555p 0.590874mV 221176.899p 0.509884mV 221186.237p 0.56202mV 221239.475p 0.385206mV 222040.799p 0.560286mV 222065.739p 0.647151mV 222086.824p 0.606853mV 223026.785p 0.620919mV 223032.012p 0.594703mV 223036.884p 0.621611mV 224013.181p 0.548085mV 224028.527p 0.465454mV 225004.164p 0.549653mV 226001.56p 0.550279mV 226031.0p 0.609255mV 226059.044p 0.699463mV 226059.763p 0.699463mV 227017.905p 0.528202mV 227074.68p 0.555238mV 227085.761p 0.474939mV 227097.897p 0.472865mV 227113.688p 0.440136mV 228003.826p 0.552858mV 228020.828p 0.548861mV 228032.389p 0.494074mV 228040.828p 0.491196mV 228059.858p 0.457329mV 229053.625p 0.538701mV 229067.153p 0.560282mV 229078.234p 0.609671mV 229093.6p 0.580569mV 229108.09p 0.607431mV 229111.668p 0.582108mV 229124.104p 0.585044mV 229124.641p 0.585044mV 229126.807p 0.560714mV 229130.469p 0.589129mV 229131.713p 0.589129mV 229144.713p 0.6463mV 230025.21p 0.474452mV 230044.863p 0.552837mV 230058.935p 0.576888mV 230060.642p 0.549714mV 230064.584p 0.549714mV 230065.994p 0.575371mV 230104.542p 0.600702mV 230109.521p 0.575599mV 230112.221p 0.550833mV 230166.445p 0.522956mV 230208.499p 0.545475mV 230214.639p 0.515116mV 230220.883p 0.454185mV 231019.392p 0.578454mV 231045.772p 0.641433mV 231046.103p 0.641433mV 231047.684p 0.641433mV 231048.393p 0.641433mV 231053.494p 0.618508mV 231062.876p 0.626464mV 232022.992p 0.44327mV 233014.42p 0.545818mV 234049.222p 0.529542mV 234059.855p 0.530516mV 234103.097p 0.505394mV 235023.996p 0.492915mV 235029.844p 0.518495mV 235040.653p 0.593657mV 235056.468p 0.669923mV 236007.962p 0.573216mV 236130.486p 0.680857mV 236140.869p 0.688139mV 237002.139p 0.552885mV 237004.701p 0.552885mV 237004.736p 0.552885mV 237005.141p 0.580377mV 237060.267p 0.525624mV 237073.102p 0.532214mV 237110.885p 0.552733mV 237123.607p 0.609676mV 237131.693p 0.562474mV 237159.049p 0.71063mV 238056.75p 0.461966mV 239006.417p 0.526479mV 239024.977p 0.60601mV 240011.17p 0.547758mV 240052.538p 0.542174mV 240068.91p 0.561386mV 240095.824p 0.545283mV 241005.4p 0.520422mV 241009.881p 0.520422mV 241011.621p 0.546954mV 241029.481p 0.573418mV 241042.075p 0.547695mV 241048.585p 0.52175mV 241058.624p 0.46965mV 241069.697p 0.521536mV 241081.521p 0.544151mV 241117.66p 0.397432mV 242011.919p 0.495943mV 242015.663p 0.469857mV 242029.599p 0.521855mV 242057.092p 0.513131mV 242097.476p 0.488332mV 242115.326p 0.573208mV 242154.478p 0.513766mV 242159.478p 0.534525mV 243021.974p 0.545642mV 243027.116p 0.518151mV 243049.587p 0.458885mV 243066.45p 0.445072mV 243067.877p 0.445072mV 244011.194p 0.496911mV 244027.47p 0.419943mV 244100.038p 0.510492mV 245031.207p 0.55517mV 245073.48p 0.627506mV 245073.771p 0.627506mV 245094.742p 0.645256mV 246003.535p 0.547328mV 246024.207p 0.603608mV 246037.208p 0.634494mV 246074.218p 0.633433mV 247003.91p 0.550549mV 247054.233p 0.617977mV 247063.568p 0.570372mV 247064.234p 0.570372mV 247072.476p 0.628683mV 248002.032p 0.55145mV 248019.652p 0.52261mV 248032.739p 0.491812mV 248035.186p 0.463567mV 248037.115p 0.463567mV 248066.023p 0.494622mV 249000.557p 0.553891mV 249001.412p 0.553891mV 249008.947p 0.580935mV 249053.642p 0.628671mV 250001.389p 0.546316mV 250009.09p 0.52108mV 250022.686p 0.550208mV 250034.17p 0.552271mV 250037.44p 0.526818mV 250041.258p 0.501379mV 250068.134p 0.529056mV 250074.303p 0.50229mV 250075.72p 0.528065mV 250146.193p 0.545011mV 250152.91p 0.51521mV 250223.348p 0.558366mV 250259.377p 0.553952mV 250260.462p 0.523228mV 251008.424p 0.52114mV 251071.314p 0.576348mV 251084.423p 0.522634mV 251121.506p 0.626743mV 251121.855p 0.626743mV 252009.035p 0.578562mV 252051.579p 0.550605mV 252067.932p 0.578437mV 253006.255p 0.57353mV 253024.884p 0.599702mV 253040.657p 0.498367mV 254018.082p 0.520507mV 254035.3p 0.57349mV 254037.602p 0.57349mV 254046.321p 0.521179mV 254046.389p 0.521179mV 254061.246p 0.547868mV 254067.784p 0.574076mV 254093.078p 0.655169mV 254100.476p 0.658992mV 254122.726p 0.673654mV 255001.567p 0.554396mV 255005.299p 0.581138mV 255009.514p 0.581138mV 255021.109p 0.609185mV 255025.337p 0.583719mV 255037.006p 0.586411mV 255058.381p 0.595525mV 256048.933p 0.638203mV 256057.483p 0.588888mV 256086.547p 0.551311mV 256169.862p 0.441981mV 257013.605p 0.498259mV 257041.2p 0.498061mV 258025.405p 0.634778mV 258039.389p 0.639178mV 258063.791p 0.579298mV 259003.23p 0.546386mV 259039.526p 0.566025mV 259054.179p 0.59033mV 259069.317p 0.562799mV 259087.415p 0.561578mV 259089.13p 0.561578mV 259127.686p 0.507924mV 259163.36p 0.477079mV 259165.651p 0.501819mV 260008.683p 0.518737mV 260021.479p 0.437128mV 260023.566p 0.437128mV 260037.007p 0.403358mV 261019.743p 0.574067mV 261039.382p 0.576978mV 261040.778p 0.551699mV 261062.197p 0.557345mV 261087.164p 0.648208mV 261088.806p 0.648208mV 261096.737p 0.604731mV 261100.592p 0.635632mV 261102.607p 0.635632mV 262012.285p 0.498306mV 262012.311p 0.498306mV 262020.901p 0.498118mV 262050.602p 0.544242mV 262059.07p 0.569583mV 262059.865p 0.569583mV 262064.013p 0.594887mV 262066.679p 0.620319mV 262081.252p 0.646309mV 262094.741p 0.648632mV 262098.527p 0.676822mV 262098.975p 0.676822mV 263027.424p 0.579233mV 263039.286p 0.526085mV 263092.109p 0.497948mV 263122.214p 0.437161mV 264058.812p 0.547559mV 264065.989p 0.500568mV 264092.663p 0.535418mV 264109.193p 0.562695mV 264113.541p 0.536378mV 264116.905p 0.510141mV 264142.216p 0.586359mV 264162.608p 0.530696mV 264167.556p 0.503662mV 265004.454p 0.553595mV 265004.936p 0.553595mV 265020.704p 0.602386mV 265051.437p 0.655784mV 265074.622p 0.614135mV 265091.66p 0.581112mV 266018.685p 0.465551mV 266049.069p 0.498572mV 267009.032p 0.575579mV 267014.617p 0.601165mV 267031.947p 0.65376mV 267042.062p 0.603845mV 267048.928p 0.632269mV 267054.163p 0.608549mV 267074.286p 0.675283mV 268000.718p 0.552087mV 268007.956p 0.579136mV 268018.65p 0.580774mV 268029.627p 0.582832mV 268056.338p 0.538126mV 268061.054p 0.513187mV 268065.693p 0.540789mV 268081.795p 0.56997mV 268091.057p 0.57158mV 268092.529p 0.57158mV 269040.52p 0.546008mV 269052.822p 0.545135mV 270012.927p 0.605445mV 270018.072p 0.631441mV 270062.795p 0.676619mV 271003.234p 0.545652mV 271006.277p 0.57295mV 271052.538p 0.614599mV 271053.491p 0.614599mV 271058.105p 0.643955mV 272023.603p 0.549262mV 272044.188p 0.547136mV 272052.471p 0.545504mV 272054.856p 0.545504mV 272063.849p 0.491446mV 272093.928p 0.478194mV 272096.798p 0.500149mV 272123.299p 0.501733mV 272131.595p 0.542926mV 272131.607p 0.542926mV 272132.15p 0.542926mV 273010.822p 0.555746mV 273013.999p 0.555746mV 273048.211p 0.531665mV 273059.807p 0.478576mV 273062.266p 0.451696mV 273102.045p 0.430943mV 274008.177p 0.57174mV 274029.199p 0.622578mV 275000.338p 0.550174mV 275012.532p 0.551135mV 275031.801p 0.659767mV 275054.308p 0.565225mV 275065.745p 0.549907mV 275070.938p 0.57944mV 275083.219p 0.586416mV 275094.028p 0.593878mV 275094.413p 0.593878mV 276022.789p 0.554535mV 276035.51p 0.58321mV 277004.477p 0.549141mV 277035.154p 0.523062mV 277039.45p 0.523062mV 277062.406p 0.489863mV 277096.592p 0.442532mV 278001.016p 0.549512mV 278018.311p 0.629094mV 278046.307p 0.589157mV 279004.218p 0.546416mV 279024.433p 0.546495mV 279056.51p 0.41049mV 279064.754p 0.433943mV 280009.141p 0.52486mV 280072.072p 0.583816mV 280087.23p 0.657654mV 280088.486p 0.657654mV 280124.947p 0.693725mV 280126.655p 0.672517mV 281003.207p 0.547601mV 281127.243p 0.586107mV 281140.234p 0.600387mV 281141.147p 0.600387mV 281191.437p 0.463382mV 281206.6p 0.528204mV 281221.943p 0.538085mV 282010.64p 0.494368mV 282013.229p 0.494368mV 282049.007p 0.506318mV 282054.293p 0.477516mV 283012.447p 0.547356mV 283012.541p 0.547356mV 283054.904p 0.661101mV 283059.394p 0.63732mV 283067.529p 0.696379mV 283070.059p 0.674784mV 284014.525p 0.546374mV 284053.697p 0.654423mV 284058.184p 0.629871mV 285002.871p 0.548111mV 285005.467p 0.52316mV 285011.079p 0.550812mV 285024.605p 0.553166mV 285026.773p 0.580515mV 285088.266p 0.661092mV 286068.634p 0.533233mV 287042.269p 0.546914mV 287048.668p 0.519421mV 288010.706p 0.544794mV 288025.477p 0.515437mV 288029.491p 0.515437mV 288033.678p 0.540547mV 288044.001p 0.590246mV 288063.605p 0.586814mV 288065.989p 0.613403mV 288077.324p 0.667423mV 288079.087p 0.667423mV 288084.033p 0.642559mV 288112.554p 0.613107mV 289003.026p 0.548119mV 289007.012p 0.574004mV 289025.29p 0.519702mV 289027.338p 0.519702mV 289031.791p 0.54516mV 289039.555p 0.570419mV 289047.699p 0.515722mV 289061.517p 0.59116mV 289066.851p 0.563668mV 289083.288p 0.587664mV 289119.593p 0.560178mV 289186.18p 0.547988mV 289197.512p 0.4916mV 289210.486p 0.510127mV 289220.743p 0.450837mV 290009.153p 0.57781mV 290034.478p 0.496272mV 290035.301p 0.468952mV 290068.893p 0.504151mV 291000.214p 0.547899mV 292028.808p 0.468429mV 292052.411p 0.43198mV 293019.926p 0.628705mV 293036.51p 0.68488mV 293037.152p 0.68488mV 293042.462p 0.713488mV 294001.338p 0.547039mV 294005.402p 0.574346mV 294016.449p 0.629068mV 294016.609p 0.629068mV 294021.433p 0.604204mV 294027.792p 0.632413mV 294029.716p 0.632413mV 294031.112p 0.660929mV 294040.065p 0.719468mV 295025.707p 0.574004mV 295026.79p 0.574004mV 295053.541p 0.708341mV 295055.227p 0.736879mV 295060.079p 0.76627mV 295062.122p 0.76627mV 295065.678p 0.744676mV 295065.849p 0.744676mV 296003.093p 0.554455mV 296006.451p 0.526812mV 296085.912p 0.482268mV 297001.002p 0.553291mV 297005.588p 0.580978mV 297031.756p 0.67006mV 298015.393p 0.528762mV 298026.181p 0.580996mV 298035.741p 0.580674mV 298044.408p 0.554297mV 298070.201p 0.553331mV 298079.797p 0.526164mV 298090.513p 0.496755mV 298095.625p 0.521258mV 298099.422p 0.521258mV 298160.763p 0.55731mV 298188.38p 0.561118mV 298201.355p 0.572793mV 298234.428p 0.598756mV 298244.572p 0.644679mV 298246.769p 0.615884mV 298252.27p 0.640156mV 298259.396p 0.664873mV 298281.959p 0.693892mV 298286.013p 0.670592mV 298286.108p 0.670592mV 298298.147p 0.6269mV 298301.66p 0.606219mV 299001.285p 0.5502mV 299073.713p 0.484573mV 299077.441p 0.455456mV 300010.491p 0.549972mV 300038.365p 0.631185mV 300057.987p 0.639299mV 300083.738p 0.579535mV 300087.656p 0.55817mV 302008.246p 0.572954mV 302042.957p 0.607526mV 302059.251p 0.641763mV 302065.108p 0.701528mV 303004.513p 0.553942mV 303019.324p 0.629885mV 303034.017p 0.550609mV 303042.564p 0.498882mV 303052.405p 0.551874mV 303068.095p 0.52492mV 303080.006p 0.548713mV 303094.032p 0.546147mV 303103.085p 0.491214mV 304018.312p 0.633475mV 304032.799p 0.715873mV 304048.768p 0.752497mV 305004.819p 0.546183mV 305012.966p 0.493111mV 305028.598p 0.516978mV 305060.088p 0.469709mV 306001.106p 0.546496mV 306010.936p 0.492465mV 306061.909p 0.589523mV 306064.225p 0.589523mV 306092.84p 0.598892mV 306100.916p 0.552313mV 306129.776p 0.436163mV 306159.4p 0.434726mV 306164.2p 0.458044mV 307005.613p 0.522432mV 307010.209p 0.548084mV 307015.852p 0.520901mV 307036.718p 0.56928mV 307077.284p 0.454249mV 307102.782p 0.466483mV 307108.566p 0.488502mV 307113.703p 0.45801mV 309034.14p 0.540678mV 309049.067p 0.56148mV 309049.882p 0.56148mV 309118.48p 0.590155mV 309184.406p 0.6236mV 309196.923p 0.660591mV 310027.457p 0.475502mV 310060.313p 0.491731mV 310070.187p 0.484995mV 310073.344p 0.484995mV 311030.266p 0.719513mV 311030.429p 0.719513mV 312018.655p 0.577407mV 312018.986p 0.577407mV 312039.429p 0.636212mV 312054.983p 0.566733mV 312079.493p 0.507672mV 312079.512p 0.507672mV 312114.765p 0.450247mV 313011.378p 0.499549mV 313027.041p 0.475976mV 313033.757p 0.502729mV 313054.812p 0.500414mV 313084.034p 0.543618mV 313086.402p 0.568121mV 313121.291p 0.638841mV 313122.248p 0.638841mV 313135.228p 0.562183mV 313160.65p 0.544399mV 313162.877p 0.544399mV 313172.192p 0.548255mV 313176.119p 0.523691mV 313186.619p 0.579529mV 313216.1p 0.697994mV 314009.469p 0.581378mV 314013.993p 0.608621mV 315003.303p 0.54803mV 315015.867p 0.465623mV 315034.721p 0.485123mV 315037.186p 0.507826mV 315053.329p 0.573788mV 315066.763p 0.587812mV 315073.159p 0.610226mV 315099.825p 0.621587mV 315108.801p 0.669745mV 315134.94p 0.697033mV 315148.53p 0.785273mV 316023.006p 0.498184mV 316042.423p 0.552482mV 316057.923p 0.525424mV 316064.0p 0.49898mV 317018.99p 0.572008mV 317026.071p 0.519787mV 317027.587p 0.519787mV 317031.912p 0.5464mV 317047.641p 0.625768mV 317073.202p 0.661322mV 317084.551p 0.722353mV 318013.996p 0.607714mV 319005.034p 0.573611mV 319006.491p 0.573611mV 319041.737p 0.555961mV 319079.747p 0.432319mV 319087.729p 0.378549mV 320011.226p 0.550463mV 320033.926p 0.498528mV 320049.132p 0.417516mV 320049.446p 0.417516mV 320060.35p 0.383454mV 321003.074p 0.55443mV 321003.63p 0.55443mV 321060.383p 0.655913mV 322008.477p 0.578678mV 322029.07p 0.636767mV 322039.122p 0.693679mV 323022.515p 0.60421mV 323023.968p 0.60421mV 323025.068p 0.578396mV 323032.965p 0.605589mV 324004.086p 0.553685mV 324056.094p 0.636552mV 324074.762p 0.613763mV 324080.474p 0.566032mV 324100.171p 0.577639mV 324109.899p 0.554468mV 324113.481p 0.583796mV 324134.779p 0.650385mV 324138.761p 0.628897mV 325034.63p 0.559275mV 325036.802p 0.534715mV 325070.492p 0.572048mV 325119.669p 0.613504mV 325159.676p 0.478609mV 325163.186p 0.506713mV 325163.336p 0.506713mV 325164.254p 0.506713mV 325167.351p 0.534399mV 325176.694p 0.53652mV 325207.702p 0.648502mV 325218.683p 0.706996mV 325221.757p 0.737159mV 326065.641p 0.640989mV 326074.39p 0.616609mV 326091.024p 0.734135mV 327002.368p 0.548991mV 327003.219p 0.548991mV 327012.058p 0.598774mV 327039.44p 0.570411mV 327040.213p 0.597619mV 327102.343p 0.440351mV 328006.387p 0.580933mV 328058.995p 0.533916mV 328091.982p 0.446256mV 329013.465p 0.492007mV 329014.574p 0.492007mV 329041.653p 0.536882mV 329057.869p 0.506477mV 329063.877p 0.478731mV 329064.394p 0.478731mV 329078.924p 0.55116mV 329104.03p 0.618103mV 329108.861p 0.590086mV 329109.972p 0.590086mV 329111.347p 0.562471mV 329112.026p 0.562471mV 329131.605p 0.612018mV 329136.547p 0.638246mV 329147.12p 0.639364mV 329160.687p 0.724585mV 330045.744p 0.636376mV 330047.236p 0.636376mV 330063.342p 0.566668mV 330081.441p 0.58159mV 330115.527p 0.533604mV 330138.181p 0.498797mV 330181.358p 0.438697mV 331033.221p 0.597328mV 331058.886p 0.683178mV 331063.869p 0.660056mV 331070.492p 0.616503mV 331080.262p 0.627071mV 331081.445p 0.627071mV 331084.42p 0.627071mV 332028.716p 0.569076mV 332033.858p 0.594715mV 332038.854p 0.620477mV 332070.922p 0.543943mV 332075.536p 0.570961mV 332125.111p 0.62992mV 332131.61p 0.657232mV 333012.992p 0.493957mV 334002.501p 0.5543mV 334034.896p 0.558332mV 334053.724p 0.508573mV 334060.638p 0.509079mV 334062.226p 0.509079mV 335005.57p 0.578192mV 335012.01p 0.60482mV 335033.118p 0.608084mV 335053.388p 0.668314mV 335063.906p 0.72789mV 336015.709p 0.633944mV 336034.303p 0.664522mV 336043.342p 0.670085mV 336044.551p 0.670085mV 336046.23p 0.700111mV 337060.323p 0.644937mV 337062.52p 0.644937mV 337073.278p 0.59281mV 337084.363p 0.542461mV 337110.007p 0.497627mV 337126.747p 0.578025mV 337174.526p 0.562031mV 337197.932p 0.652265mV 337213.182p 0.585305mV 338014.731p 0.495889mV 338036.079p 0.627129mV 338045.688p 0.575364mV 338055.447p 0.524926mV 338056.827p 0.524926mV 338058.433p 0.524926mV 338078.479p 0.582018mV 338079.353p 0.582018mV 338143.682p 0.632054mV 338146.538p 0.609585mV 339000.285p 0.547431mV 339019.325p 0.51891mV 339058.994p 0.50218mV 339063.95p 0.472668mV 340055.668p 0.736931mV 341044.365p 0.442977mV 341051.107p 0.49244mV 341067.074p 0.458119mV 341068.749p 0.458119mV 341069.912p 0.458119mV 342023.74p 0.489574mV 343005.585p 0.520235mV 343025.736p 0.628422mV 343027.112p 0.628422mV 343029.397p 0.628422mV 343050.986p 0.558772mV 343092.811p 0.52519mV 343121.105p 0.693457mV 343121.931p 0.693457mV 343125.54p 0.670542mV 343125.97p 0.670542mV 344048.697p 0.585524mV 344075.918p 0.486681mV 344106.142p 0.42717mV 346031.891p 0.450924mV 346041.801p 0.50334mV 346048.3p 0.476113mV 346050.302p 0.448607mV 346080.427p 0.484367mV 347043.95p 0.596836mV 347048.405p 0.570131mV 347069.522p 0.46458mV 347088.161p 0.45983mV 347099.923p 0.455079mV 347118.645p 0.438288mV 348088.605p 0.510407mV 348089.014p 0.510407mV 349024.912p 0.442561mV 349030.293p 0.438953mV 350016.477p 0.52218mV 350032.805p 0.54742mV 350103.681p 0.514541mV 350106.1p 0.483417mV 350109.114p 0.483417mV 351027.419p 0.479525mV 352019.503p 0.519419mV 352027.544p 0.569912mV 352043.852p 0.540192mV 352048.228p 0.512539mV 352059.356p 0.509503mV 352094.559p 0.568855mV 352132.027p 0.650612mV 352144.836p 0.648057mV 352160.527p 0.649957mV 353009.71p 0.519657mV 353031.962p 0.536567mV 353060.611p 0.516587mV 353082.187p 0.603144mV 353093.364p 0.543027mV 353163.752p 0.535068mV 354000.511p 0.548549mV 354012.972p 0.54617mV 354031.93p 0.540155mV 354057.948p 0.610301mV 354066.946p 0.607449mV 354088.028p 0.606509mV 354090.983p 0.633253mV 354103.323p 0.635276mV 354108.227p 0.66321mV 354132.233p 0.601652mV 354135.822p 0.580668mV 355046.384p 0.535524mV 355048.703p 0.535524mV 355069.422p 0.591512mV 355104.153p 0.579767mV 355108.234p 0.55668mV 355132.871p 0.546821mV 355139.484p 0.523674mV 355147.713p 0.581877mV 355160.534p 0.669676mV 356011.887p 0.550507mV 356032.058p 0.547259mV 356041.762p 0.546078mV 356048.092p 0.518961mV 357032.179p 0.597776mV 357035.236p 0.623969mV 357037.302p 0.623969mV 357081.946p 0.770855mV 358037.554p 0.680522mV 358040.051p 0.708125mV 358046.561p 0.736479mV 359019.328p 0.576916mV 359039.739p 0.576544mV 359049.543p 0.629545mV 359051.924p 0.656456mV 359059.589p 0.683848mV 359084.649p 0.673995mV 361010.687p 0.597841mV 361020.129p 0.597726mV 361028.036p 0.624294mV 361069.472p 0.64507mV 362001.034p 0.552032mV 362048.989p 0.647365mV 362054.978p 0.677348mV 363034.203p 0.498546mV 363079.351p 0.521732mV 363101.812p 0.59653mV 363119.946p 0.568851mV 363164.634p 0.502219mV 363185.863p 0.430113mV 363192.994p 0.455999mV 364025.634p 0.524832mV 364052.387p 0.655236mV 364055.017p 0.682144mV 364058.6p 0.682144mV 365060.049p 0.602973mV 365120.453p 0.683031mV 366008.062p 0.523141mV 366050.52p 0.579972mV 366103.261p 0.724074mV 366104.641p 0.724074mV 366108.367p 0.700043mV 366117.033p 0.707451mV 366118.318p 0.707451mV 367000.397p 0.553885mV 367020.162p 0.498148mV 367020.239p 0.498148mV 367020.366p 0.498148mV 367034.398p 0.547286mV 367039.017p 0.518972mV 367076.231p 0.603178mV 367088.695p 0.547404mV 367099.797p 0.59747mV 367122.21p 0.674353mV 368027.323p 0.520024mV 368028.306p 0.520024mV 368066.236p 0.560577mV 368073.55p 0.533458mV 368086.35p 0.504812mV 368090.619p 0.530256mV 368095.638p 0.502772mV 368116.28p 0.495011mV 368151.766p 0.443193mV 369019.984p 0.57768mV 369039.812p 0.687414mV 369050.111p 0.722939mV 370009.487p 0.525988mV 370013.109p 0.498931mV 370020.548p 0.49687mV 370048.956p 0.566075mV 370051.145p 0.589829mV 370097.395p 0.665664mV 370097.487p 0.665664mV 370106.602p 0.672846mV 370112.928p 0.703543mV 371005.085p 0.520138mV 371032.062p 0.487597mV 371059.463p 0.503821mV 371065.279p 0.445434mV 371077.548p 0.43746mV 372014.698p 0.543343mV 372031.073p 0.589941mV 372062.36p 0.531997mV 372075.36p 0.450789mV 372086.533p 0.394786mV 373027.215p 0.572549mV 373043.513p 0.60003mV 373046.375p 0.574255mV 373055.86p 0.628808mV 373073.939p 0.607903mV 373087.59p 0.643507mV 373089.525p 0.643507mV 373098.924p 0.652608mV 374012.465p 0.60699mV 374033.995p 0.614648mV 374052.995p 0.627216mV 374078.512p 0.521166mV 374082.653p 0.500395mV 374094.25p 0.458051mV 374111.143p 0.471765mV 374115.723p 0.500622mV 374118.417p 0.500622mV 374132.252p 0.427185mV 375012.143p 0.551811mV 375025.256p 0.527004mV 375034.846p 0.553443mV 376023.708p 0.600434mV 376042.002p 0.549296mV 376074.39p 0.559088mV 376079.093p 0.587973mV 376092.442p 0.62288mV 377001.453p 0.550193mV 377018.459p 0.520517mV 377033.843p 0.541313mV 377072.426p 0.569385mV 377087.69p 0.636497mV 377106.727p 0.680408mV 377107.079p 0.680408mV 377118.959p 0.68049mV 377143.982p 0.720848mV 378009.396p 0.519445mV 378013.989p 0.492737mV 378048.839p 0.509793mV 378061.505p 0.527236mV 378150.319p 0.583048mV 378180.045p 0.624015mV 378192.697p 0.622735mV 378193.882p 0.622735mV 378194.873p 0.622735mV 378208.282p 0.651261mV 378222.168p 0.631981mV 378237.309p 0.669528mV 378239.591p 0.669528mV 379004.197p 0.549194mV 379076.157p 0.552797mV 379094.314p 0.5682mV 379098.148p 0.538896mV 379114.371p 0.503566mV 380003.366p 0.552414mV 380021.113p 0.557704mV 380033.469p 0.50847mV 380065.823p 0.540562mV 380066.138p 0.540562mV 380101.872p 0.515651mV 380106.832p 0.489811mV 380125.541p 0.488998mV 380154.088p 0.507139mV 380189.891p 0.613505mV 380206.176p 0.65498mV 380209.895p 0.65498mV 380311.732p 0.548187mV 380317.787p 0.574789mV 380344.505p 0.496943mV 380349.795p 0.470327mV 380368.583p 0.464496mV 381006.517p 0.522572mV 381029.482p 0.464703mV 381035.931p 0.460077mV 381042.044p 0.482949mV 381050.42p 0.526922mV 382000.427p 0.550229mV 382025.327p 0.583496mV 382043.199p 0.668618mV 382059.934p 0.653424mV 383028.152p 0.624407mV 383076.742p 0.74598mV 384023.234p 0.599644mV 384036.823p 0.679651mV 384036.972p 0.679651mV 384039.463p 0.679651mV 384039.951p 0.679651mV 384058.68p 0.743057mV 385013.369p 0.498343mV 385027.718p 0.471953mV 386000.336p 0.549392mV 386007.231p 0.574966mV 386027.979p 0.519529mV 386031.138p 0.545038mV 386042.023p 0.542982mV 386063.928p 0.589958mV 386080.186p 0.638837mV 386105.882p 0.511946mV 386113.545p 0.539584mV 387061.535p 0.611081mV 387065.102p 0.640564mV 387070.076p 0.670367mV 388020.393p 0.599389mV 388027.579p 0.573253mV 388079.133p 0.641887mV 388111.72p 0.538284mV 388126.944p 0.523829mV 388134.72p 0.553778mV 388155.969p 0.65258mV 389020.799p 0.496156mV 389021.011p 0.496156mV 389040.397p 0.48634mV 389061.707p 0.522286mV 390014.318p 0.553281mV 390019.181p 0.52724mV 390033.042p 0.554273mV 391011.745p 0.551272mV 391029.475p 0.579663mV 391036.832p 0.634779mV 391048.087p 0.638662mV 391065.155p 0.651614mV 391066.178p 0.651614mV 392030.572p 0.548858mV 392031.256p 0.548858mV 392034.309p 0.548858mV 393028.843p 0.52746mV 393033.409p 0.500899mV 393081.384p 0.43257mV 394016.259p 0.517823mV 394028.531p 0.515292mV 394031.892p 0.539838mV 394035.394p 0.511611mV 394035.453p 0.511611mV 395018.113p 0.468203mV 395023.607p 0.493324mV 395024.508p 0.493324mV 396000.827p 0.552903mV 396011.442p 0.554339mV 396031.002p 0.61148mV 396071.667p 0.685187mV 396078.037p 0.663725mV 397019.924p 0.523949mV 397056.561p 0.40597mV 398006.901p 0.572709mV 398032.076p 0.600543mV 398045.008p 0.526858mV 398060.627p 0.558411mV 398071.526p 0.561224mV 398090.757p 0.62158mV 398094.279p 0.62158mV 398096.723p 0.650741mV 398107.933p 0.606076mV 398111.022p 0.584674mV 398139.204p 0.58442mV 399004.314p 0.549001mV 399031.759p 0.494862mV 399045.808p 0.516588mV 399063.554p 0.482509mV 400041.896p 0.565693mV 400046.27p 0.540995mV 400066.449p 0.546856mV 400110.286p 0.416082mV 400144.76p 0.445862mV 401019.241p 0.524905mV 401027.811p 0.575996mV 401060.645p 0.488344mV 401064.083p 0.488344mV 401093.458p 0.571734mV 401102.976p 0.564247mV 401119.134p 0.528303mV 401123.0p 0.551446mV 402002.885p 0.553222mV 402047.347p 0.582452mV 402071.275p 0.560781mV 402146.624p 0.567885mV 402147.497p 0.567885mV 402161.432p 0.549369mV 402161.646p 0.549369mV 402168.18p 0.578mV 402187.141p 0.694049mV 403000.607p 0.554383mV 403051.071p 0.554493mV 403101.67p 0.598753mV 403126.493p 0.526378mV 403132.93p 0.554238mV 403135.275p 0.529349mV 403139.016p 0.529349mV 403167.939p 0.591839mV 403185.564p 0.60425mV 403191.087p 0.581941mV 403195.638p 0.612071mV 404004.546p 0.549012mV 404014.743p 0.604168mV 404016.786p 0.579294mV 404023.92p 0.607348mV 404054.835p 0.625816mV 405041.666p 0.506217mV 405045.135p 0.480653mV 405062.052p 0.506992mV 406012.869p 0.602854mV 406041.443p 0.613879mV 406095.733p 0.469203mV 406098.109p 0.469203mV 406101.46p 0.498089mV 406146.378p 0.481857mV 406175.595p 0.577838mV 406224.441p 0.477933mV 406233.039p 0.418371mV 407001.467p 0.546992mV 407011.526p 0.596889mV 407022.188p 0.594718mV 407034.508p 0.594044mV 407083.933p 0.610426mV 407087.781p 0.587757mV 407095.526p 0.595677mV 407104.035p 0.62612mV 408011.531p 0.601732mV 408019.987p 0.574569mV 408022.167p 0.547723mV 408027.851p 0.573708mV 408059.959p 0.57271mV 408074.455p 0.547998mV 408076.663p 0.575265mV 408116.675p 0.529878mV 408117.374p 0.529878mV 408130.153p 0.505483mV 408151.603p 0.505201mV 408176.227p 0.470033mV 408176.768p 0.470033mV 409006.264p 0.579828mV 409011.033p 0.606877mV 409020.877p 0.661678mV 409022.919p 0.661678mV 409028.968p 0.68974mV 409034.4p 0.718433mV 409039.352p 0.747877mV 410000.044p 0.550606mV 410004.144p 0.550606mV 410010.911p 0.500326mV 410023.761p 0.502066mV 410024.576p 0.502066mV 410056.597p 0.468902mV 410060.507p 0.439957mV 411013.398p 0.605872mV 411018.727p 0.580955mV 411029.157p 0.584644mV 411039.252p 0.589491mV 412012.759p 0.544164mV 412028.999p 0.567806mV 412029.483p 0.567806mV 412039.034p 0.513511mV 412044.591p 0.486362mV 412061.395p 0.533007mV 412061.509p 0.533007mV 412062.659p 0.533007mV 412074.297p 0.476304mV 413042.683p 0.584735mV 413046.643p 0.609632mV 413071.738p 0.527724mV 413073.851p 0.527724mV 413076.354p 0.501356mV 413085.697p 0.448038mV 413091.666p 0.47342mV 413091.752p 0.47342mV 413102.946p 0.469799mV 413110.17p 0.516931mV 413119.944p 0.539822mV 413127.566p 0.585062mV 413195.595p 0.6196mV 413219.568p 0.625497mV 413225.987p 0.683117mV 413229.007p 0.683117mV 413237.349p 0.690964mV 413237.814p 0.690964mV 414015.365p 0.58309mV 414032.812p 0.510458mV 414035.514p 0.538779mV 414045.206p 0.542328mV 414068.033p 0.548857mV 414120.581p 0.518706mV 414172.232p 0.538883mV 414173.902p 0.538883mV 414175.767p 0.509106mV 414177.943p 0.509106mV 414181.131p 0.479273mV 414184.238p 0.479273mV 414196.947p 0.387951mV 415001.074p 0.552357mV 415004.473p 0.552357mV 416058.903p 0.551336mV 416072.848p 0.591765mV 416088.363p 0.581475mV 417028.297p 0.587686mV 417037.528p 0.643688mV 417053.277p 0.678473mV 418005.47p 0.521934mV 418021.308p 0.54423mV 418075.444p 0.495514mV 418087.175p 0.488935mV 418094.461p 0.458929mV 418103.964p 0.449628mV 419021.008p 0.555141mV 419025.351p 0.582173mV 419051.779p 0.668546mV 419053.151p 0.668546mV 420005.712p 0.522207mV 420017.728p 0.575844mV 420020.572p 0.549894mV 420038.078p 0.578047mV 420116.968p 0.414111mV 421001.075p 0.552218mV 421006.189p 0.579021mV 421023.37p 0.607522mV 421068.492p 0.604414mV 421081.024p 0.591026mV 421087.949p 0.62152mV 421096.059p 0.579811mV 421100.111p 0.559602mV 422009.437p 0.575656mV 422023.38p 0.495725mV 422060.804p 0.429086mV 422066.244p 0.39907mV 423001.47p 0.553179mV 423002.839p 0.553179mV 423023.727p 0.495076mV 423024.666p 0.495076mV 423060.245p 0.528566mV 423092.146p 0.615883mV 423109.969p 0.585686mV 423124.956p 0.557033mV 423125.015p 0.529919mV 423129.043p 0.529919mV 425085.905p 0.552746mV 425098.1p 0.553145mV 425119.265p 0.553176mV 425144.416p 0.632785mV 426005.924p 0.576583mV 426057.476p 0.540346mV 426071.194p 0.622945mV 426074.184p 0.622945mV 426080.413p 0.67907mV 426087.089p 0.655488mV 427002.384p 0.550983mV 427004.452p 0.550983mV 427010.404p 0.551087mV 427012.68p 0.551087mV 427028.049p 0.629983mV 427040.022p 0.659196mV 427040.758p 0.659196mV 428006.027p 0.524063mV 428016.302p 0.52349mV 428024.621p 0.549124mV 428026.848p 0.521931mV 428064.666p 0.647365mV 428065.565p 0.620945mV 428078.687p 0.622446mV 428100.19p 0.658868mV 428114.166p 0.666044mV 429001.596p 0.550933mV 429003.079p 0.550933mV 429006.804p 0.576579mV 429016.794p 0.575383mV 429037.155p 0.574941mV 429042.902p 0.548389mV 429060.016p 0.442089mV 430004.559p 0.548975mV 430004.59p 0.548975mV 430004.985p 0.548975mV 431038.626p 0.518823mV 431044.464p 0.493093mV 431070.751p 0.488774mV 432051.632p 0.620559mV 432073.727p 0.688692mV 433041.896p 0.481889mV 433084.485p 0.500505mV 434001.139p 0.547345mV 434008.699p 0.520275mV 434010.754p 0.493189mV 434012.886p 0.493189mV 435005.373p 0.51962mV 435015.864p 0.517966mV 435017.055p 0.517966mV 435047.448p 0.453177mV 435047.897p 0.453177mV 435063.214p 0.466319mV 436066.529p 0.557575mV 436068.306p 0.557575mV 436100.138p 0.678306mV 437011.353p 0.554378mV 437033.819p 0.451446mV 437046.826p 0.475668mV 437048.85p 0.475668mV 437067.062p 0.465081mV 437068.271p 0.465081mV 438012.549p 0.547229mV 438034.306p 0.594085mV 438055.795p 0.509766mV 438071.478p 0.530211mV 439043.67p 0.546776mV 439048.266p 0.573414mV 439127.297p 0.54335mV 439142.577p 0.470429mV 439156.153p 0.447154mV 439176.009p 0.390555mV 439187.689p 0.434884mV 440015.69p 0.570286mV 440025.065p 0.516031mV 440039.14p 0.46161mV 440045.059p 0.510888mV 440062.856p 0.476793mV 440067.375p 0.499666mV 440068.372p 0.499666mV 440072.343p 0.469858mV 440091.608p 0.503212mV 441001.061p 0.55295mV 441011.592p 0.603499mV 441035.169p 0.628545mV 441041.082p 0.655665mV 441053.618p 0.658917mV 441057.596p 0.687883mV 441062.309p 0.665201mV 441074.377p 0.674386mV 442007.147p 0.526591mV 442010.89p 0.5533mV 442015.885p 0.579863mV 442018.018p 0.579863mV 442035.898p 0.635287mV 442042.083p 0.663245mV 442046.125p 0.63919mV 442056.788p 0.645618mV 442063.389p 0.675819mV 443070.086p 0.463363mV 443097.486p 0.481796mV 443132.659p 0.480116mV 444034.964p 0.537089mV 444056.449p 0.663696mV 444093.04p 0.542059mV 444096.851p 0.570642mV 444102.692p 0.546692mV 444122.671p 0.50317mV 445023.07p 0.499196mV 445071.208p 0.376048mV 446038.644p 0.466108mV 447005.303p 0.580298mV 447016.591p 0.634408mV 447026.666p 0.689888mV 447027.869p 0.689888mV 447032.369p 0.666045mV 447046.669p 0.599772mV 447051.573p 0.578936mV 447052.955p 0.578936mV 448001.896p 0.547458mV 448003.021p 0.547458mV 448038.635p 0.463288mV 449003.161p 0.54735mV 449004.104p 0.54735mV 449013.872p 0.549364mV 449019.147p 0.576836mV 449042.891p 0.504781mV 449051.218p 0.507307mV 449058.964p 0.534646mV 449061.373p 0.509063mV 449084.754p 0.456796mV 449109.178p 0.524523mV 449127.256p 0.512806mV 449147.441p 0.444643mV 450008.112p 0.573316mV 450037.112p 0.68663mV 450049.755p 0.745253mV 451017.09p 0.521862mV 451030.817p 0.546225mV 452000.084p 0.549373mV 452004.924p 0.549373mV 452007.917p 0.522172mV 452128.218p 0.688992mV 453021.416p 0.557175mV 453028.505p 0.532451mV 453094.326p 0.560666mV 453109.261p 0.584811mV 453118.031p 0.584706mV 453124.993p 0.558475mV 453158.909p 0.480454mV 454002.215p 0.551315mV 455002.369p 0.551291mV 455050.965p 0.485828mV 455054.023p 0.485828mV 455072.335p 0.424134mV 456005.529p 0.522803mV 456016.143p 0.47076mV 456043.69p 0.440296mV 457002.548p 0.548174mV 457003.156p 0.548174mV 457007.901p 0.521534mV 457015.407p 0.468055mV 457029.841p 0.465852mV 458020.875p 0.555654mV 458024.469p 0.555654mV 458058.04p 0.646222mV 458062.684p 0.675381mV 458068.994p 0.70505mV 459007.232p 0.526236mV 459012.36p 0.551711mV 460024.657p 0.655468mV 460031.987p 0.603803mV 460036.0p 0.631446mV 460040.158p 0.659404mV 460050.506p 0.716857mV 461019.26p 0.529903mV 461066.644p 0.656221mV 462000.871p 0.551723mV 462009.64p 0.52494mV 462010.725p 0.550843mV 462011.872p 0.550843mV 462023.514p 0.549663mV 464006.491p 0.52528mV 464009.226p 0.52528mV 464034.659p 0.494604mV 464057.914p 0.511018mV 464086.301p 0.486485mV 465005.652p 0.5276mV 466021.679p 0.490482mV 466032.93p 0.487386mV 466049.909p 0.400644mV 467037.184p 0.520498mV 468015.534p 0.527802mV 468032.796p 0.450165mV 468037.993p 0.423572mV 468065.367p 0.458503mV 470006.592p 0.574021mV 470007.102p 0.574021mV 470019.125p 0.574785mV 470022.244p 0.549231mV 470065.218p 0.478969mV 470113.093p 0.497307mV 470128.601p 0.460222mV 471036.659p 0.519165mV 471054.656p 0.434545mV 471055.937p 0.405573mV 471063.356p 0.428202mV 471073.448p 0.470486mV 472003.214p 0.551847mV 472018.41p 0.632351mV 472048.574p 0.644955mV 472064.058p 0.632238mV 473006.017p 0.574398mV 473015.178p 0.576542mV 473017.633p 0.576542mV 473048.832p 0.587075mV 473059.43p 0.644656mV 473061.107p 0.621586mV 473079.07p 0.71213mV 474007.537p 0.523963mV 474053.098p 0.382091mV 475009.573p 0.579254mV 475033.474p 0.609672mV 475038.6p 0.637007mV 475039.353p 0.637007mV 475042.05p 0.612086mV 475044.979p 0.612086mV 475049.142p 0.587749mV 475053.594p 0.563836mV 475078.485p 0.65796mV 476040.64p 0.555367mV 476106.493p 0.605875mV 477005.104p 0.577051mV 477009.856p 0.577051mV 477026.088p 0.631304mV 477036.808p 0.581011mV 477054.501p 0.665884mV 477066.668p 0.650415mV 478005.675p 0.575784mV 478008.778p 0.575784mV 478008.953p 0.575784mV 478036.589p 0.526588mV 478069.803p 0.530229mV 478071.025p 0.503539mV 479010.395p 0.548496mV 479023.377p 0.545559mV 479044.36p 0.539056mV 479049.188p 0.511257mV 479050.604p 0.483393mV 479071.284p 0.420932mV 480018.818p 0.519787mV 480021.785p 0.545726mV 480023.554p 0.545726mV 480036.9p 0.517366mV 481003.723p 0.545941mV 481011.773p 0.548279mV 481045.904p 0.478035mV 481064.674p 0.451904mV 481077.943p 0.472685mV 481083.094p 0.443534mV 481096.066p 0.456837mV 482004.539p 0.551472mV 482030.15p 0.59823mV 482076.042p 0.641682mV 483033.542p 0.609238mV 484045.516p 0.58895mV 484063.501p 0.568849mV 484128.559p 0.579017mV 484139.884p 0.587595mV 484140.153p 0.566061mV 484156.971p 0.554716mV 484175.505p 0.62773mV 484179.529p 0.62773mV 485040.25p 0.553262mV 485074.545p 0.555321mV 485139.61p 0.434761mV 485158.589p 0.428611mV 485170.963p 0.441915mV 486003.341p 0.548263mV 486019.579p 0.519053mV 486031.486p 0.488632mV 486061.609p 0.467213mV 487027.02p 0.631085mV 487038.455p 0.635104mV 487061.725p 0.681335mV 488006.038p 0.580372mV 488007.282p 0.580372mV 488029.419p 0.528033mV 488033.538p 0.502009mV 488039.731p 0.475844mV 488092.931p 0.428813mV 488103.444p 0.367896mV 489033.729p 0.552543mV 489080.708p 0.502525mV 489123.691p 0.610914mV 489151.901p 0.565376mV 489156.491p 0.540697mV 489170.421p 0.624687mV 489174.797p 0.624687mV 489191.397p 0.582667mV 489192.447p 0.582667mV 489195.521p 0.612159mV 489202.73p 0.641822mV 490001.204p 0.547885mV 490001.73p 0.547885mV 490030.956p 0.500378mV 490056.425p 0.524373mV 490062.464p 0.550009mV 490083.622p 0.598865mV 490107.544p 0.678116mV 490119.872p 0.735815mV 491039.478p 0.465165mV 491067.837p 0.444495mV 492031.53p 0.442966mV 493075.953p 0.611543mV 493082.348p 0.59088mV 494020.988p 0.550629mV 494027.846p 0.5252mV 494043.235p 0.553931mV 494050.333p 0.607851mV 494052.803p 0.607851mV 494056.028p 0.635012mV 494066.002p 0.690526mV 494081.448p 0.726866mV 495022.171p 0.544644mV 495032.202p 0.541126mV 495033.591p 0.541126mV 495039.66p 0.51318mV 495044.389p 0.537755mV 495049.019p 0.509541mV 495058.969p 0.557756mV 495080.041p 0.572103mV 495083.859p 0.572103mV 495085.485p 0.59642mV 495091.016p 0.568328mV 495141.933p 0.391589mV 496019.715p 0.5259mV 496035.292p 0.476337mV 496048.699p 0.423545mV 496079.93p 0.459198mV 497005.148p 0.527681mV 497007.454p 0.527681mV 497017.56p 0.526694mV 497017.755p 0.526694mV 497030.146p 0.498132mV 497062.323p 0.48816mV 497068.256p 0.511968mV 497074.079p 0.535347mV 497077.65p 0.55846mV 497079.316p 0.55846mV 497085.878p 0.499905mV 497150.938p 0.577906mV 497159.803p 0.548149mV 497177.199p 0.63918mV 497189.325p 0.581909mV 497194.084p 0.606439mV 497195.523p 0.578593mV 497203.667p 0.60371mV 497220.273p 0.601975mV 497257.901p 0.582357mV 497264.057p 0.610797mV 497279.682p 0.645091mV 497298.527p 0.661417mV 498043.769p 0.536304mV 498085.512p 0.53948mV 498120.572p 0.441844mV 499001.966p 0.552451mV 500028.575p 0.631327mV 500029.639p 0.631327mV 500036.628p 0.635195mV 500043.464p 0.663972mV 501029.265p 0.480766mV 501033.728p 0.507387mV 502019.985p 0.574469mV 502064.802p 0.554891mV 502079.087p 0.635871mV 502108.502p 0.596272mV 503004.366p 0.549224mV 504007.493p 0.580201mV 504021.936p 0.555788mV 504023.181p 0.555788mV 504061.998p 0.509101mV 505002.572p 0.548457mV 505004.36p 0.548457mV 505014.637p 0.495974mV 505046.862p 0.455862mV 506000.959p 0.545681mV 506012.654p 0.54643mV 506038.577p 0.468374mV 506054.119p 0.492176mV 506056.251p 0.516467mV 506104.435p 0.509598mV 507019.152p 0.581129mV 507026.266p 0.584142mV 507027.411p 0.584142mV 507034.569p 0.559501mV 507040.936p 0.510742mV 507058.855p 0.48907mV 507060.413p 0.46336mV 508021.909p 0.65546mV 508026.234p 0.681856mV 508036.298p 0.684076mV 508050.273p 0.667372mV 509013.368p 0.497414mV 509062.979p 0.709573mV 509063.837p 0.709573mV 510039.089p 0.568817mV 510050.966p 0.591155mV 510068.739p 0.563762mV 510104.669p 0.542415mV 510113.564p 0.491957mV 510138.22p 0.571326mV 510167.869p 0.569282mV 510174.384p 0.595939mV 510192.51p 0.546111mV 510193.959p 0.546111mV 510216.41p 0.46934mV 510232.323p 0.441282mV 511026.691p 0.571933mV 511035.562p 0.570624mV 511039.073p 0.570624mV 511062.885p 0.650817mV 511065.212p 0.678474mV 512003.834p 0.547561mV 512082.903p 0.479403mV 512090.645p 0.523313mV 512117.398p 0.525858mV 512117.889p 0.525858mV 512118.912p 0.525858mV 512140.243p 0.581436mV 512196.306p 0.575518mV 512209.093p 0.573564mV 512219.361p 0.571894mV 512224.781p 0.544778mV 512257.023p 0.562089mV 512262.362p 0.586181mV 512267.657p 0.610357mV 512290.275p 0.683443mV 512303.741p 0.684848mV 512306.562p 0.660698mV 512309.621p 0.660698mV 512309.826p 0.660698mV 513029.439p 0.582735mV 513033.614p 0.557636mV 513037.012p 0.58536mV 513052.393p 0.669444mV 513053.878p 0.669444mV 514035.76p 0.468507mV 515005.602p 0.575072mV 515015.913p 0.626374mV 515060.719p 0.61699mV 516020.209p 0.493512mV 516062.828p 0.472902mV 516074.119p 0.517774mV 516089.286p 0.530607mV 516100.322p 0.542634mV 516161.037p 0.53503mV 516161.598p 0.53503mV 516188.902p 0.537338mV 517001.255p 0.550824mV 517032.253p 0.604297mV 517046.822p 0.687341mV 519037.32p 0.474982mV 519047.328p 0.526845mV 519047.855p 0.526845mV 519098.049p 0.50977mV 520020.745p 0.545313mV 520065.522p 0.506647mV 520083.89p 0.474313mV 520102.738p 0.566713mV 520116.058p 0.477947mV 521018.001p 0.523016mV 521020.928p 0.548959mV 521025.875p 0.522059mV 521037.782p 0.520736mV 521045.835p 0.518359mV 522021.505p 0.49605mV 522028.55p 0.469535mV 522052.813p 0.435878mV 523038.139p 0.573297mV 523075.353p 0.454023mV 524016.711p 0.627666mV 524020.794p 0.655237mV 524038.72p 0.741228mV 525008.205p 0.519636mV 525019.731p 0.572892mV 525027.34p 0.626055mV 525027.746p 0.626055mV 525038.877p 0.627767mV 525055.95p 0.689665mV 525062.795p 0.720011mV 526007.401p 0.576396mV 526058.89p 0.529467mV 526063.64p 0.503831mV 526072.178p 0.504676mV 526078.031p 0.530838mV 527008.493p 0.578936mV 527020.104p 0.656383mV 527023.007p 0.656383mV 527035.596p 0.685737mV 528017.181p 0.575456mV 528023.485p 0.549797mV 528058.944p 0.529999mV 528059.273p 0.529999mV 528060.286p 0.557732mV 528067.171p 0.585345mV 528067.982p 0.585345mV 528071.468p 0.613003mV 528111.328p 0.524365mV 528142.898p 0.427375mV 528177.861p 0.440208mV 529002.822p 0.547413mV 529034.955p 0.603104mV 529054.251p 0.662237mV 530011.098p 0.606122mV 530021.461p 0.556041mV 531021.441p 0.547125mV 531082.935p 0.598413mV 532002.233p 0.55155mV 532063.557p 0.526118mV 532070.408p 0.568677mV 532098.807p 0.520898mV 532105.986p 0.565221mV 532127.392p 0.60135mV 532149.064p 0.588462mV 532212.647p 0.731074mV 533006.783p 0.527281mV 533041.703p 0.604468mV 533087.596p 0.415983mV 534009.37p 0.57227mV 534020.598p 0.595732mV 534039.98p 0.621352mV 534042.043p 0.648129mV 534051.911p 0.703135mV 534052.96p 0.703135mV 534064.045p 0.760982mV 534064.867p 0.760982mV 535009.038p 0.521787mV 535015.228p 0.521578mV 535056.393p 0.517782mV 535079.121p 0.565958mV 535088.64p 0.615537mV 535091.934p 0.588022mV 535125.115p 0.667886mV 536007.679p 0.57946mV 536014.196p 0.552837mV 536035.781p 0.525522mV 536056.014p 0.522866mV 536061.97p 0.548206mV 536089.533p 0.516267mV 536115.98p 0.452412mV 537040.243p 0.496293mV 537045.737p 0.522067mV 537071.242p 0.490748mV 538035.374p 0.472374mV 538045.687p 0.524603mV 538048.93p 0.524603mV 538050.277p 0.49748mV 539000.582p 0.545823mV 539055.363p 0.511752mV 539057.16p 0.511752mV 540011.459p 0.543717mV 540018.755p 0.568489mV 540037.051p 0.563509mV 540076.96p 0.559816mV 540140.858p 0.469093mV 541006.043p 0.524132mV 541014.802p 0.549343mV 541038.816p 0.516895mV 541071.761p 0.475262mV 541075.021p 0.498186mV 541081.626p 0.520578mV 541098.866p 0.482139mV 542031.451p 0.502863mV 542038.776p 0.530191mV 542048.199p 0.58415mV 542074.781p 0.615131mV 542093.155p 0.676435mV 542096.644p 0.706255mV 542097.97p 0.706255mV 543064.128p 0.592798mV 543108.635p 0.584255mV 543159.115p 0.464988mV 543206.616p 0.405878mV 543206.871p 0.405878mV 544002.756p 0.551005mV 544053.074p 0.539182mV 544055.761p 0.511667mV 544077.099p 0.558026mV 544104.965p 0.521046mV 544105.077p 0.492332mV 544107.405p 0.492332mV 545007.15p 0.519677mV 545030.484p 0.544205mV 545074.287p 0.53688mV 545100.871p 0.423131mV 546020.246p 0.66083mV 546028.362p 0.635691mV 546053.755p 0.677255mV 547020.852p 0.600873mV 547045.414p 0.680112mV 547049.6p 0.680112mV 547058.114p 0.736473mV 547068.022p 0.744291mV 548001.365p 0.546314mV 548023.156p 0.497292mV 548034.13p 0.49855mV 548047.02p 0.523638mV 548052.158p 0.548779mV 548056.877p 0.573745mV 548063.468p 0.598703mV 548065.732p 0.623819mV 548088.359p 0.569696mV 548132.952p 0.661772mV 549005.052p 0.528779mV 549018.081p 0.530255mV 549042.336p 0.560622mV 549049.873p 0.535779mV 549086.646p 0.488656mV 549088.696p 0.488656mV 550036.568p 0.625106mV 550049.352p 0.678099mV 550051.038p 0.705445mV 551005.681p 0.522692mV 551021.325p 0.603176mV 551032.119p 0.604699mV 552011.651p 0.549587mV 552028.864p 0.575514mV 552044.148p 0.656059mV 553009.117p 0.579836mV 553046.9p 0.523979mV 553051.294p 0.54966mV 553058.287p 0.522514mV 553079.255p 0.465879mV 554026.08p 0.41874mV 554046.566p 0.409744mV 554051.633p 0.379102mV 555028.166p 0.636095mV 556015.834p 0.525313mV 556021.771p 0.551424mV 556026.175p 0.577377mV 556035.022p 0.576796mV 556042.349p 0.60327mV 556042.967p 0.60327mV 556049.82p 0.629911mV 556073.482p 0.665877mV 556081.646p 0.675049mV 557016.41p 0.572849mV 557018.495p 0.572849mV 557019.904p 0.572849mV 557052.664p 0.598872mV 557065.871p 0.679922mV 557079.55p 0.736696mV 557080.987p 0.766288mV 558000.143p 0.550428mV 558057.133p 0.578825mV 558073.454p 0.664041mV 558074.39p 0.664041mV 558078.469p 0.640836mV 558085.89p 0.700837mV 559003.526p 0.552106mV 559011.864p 0.55314mV 559018.375p 0.579853mV 559047.214p 0.582774mV 559073.494p 0.506575mV 559098.7p 0.426592mV 559119.294p 0.468918mV 560006.645p 0.573583mV 560025.744p 0.570658mV 560025.881p 0.570658mV 560029.89p 0.570658mV 560034.237p 0.597115mV 560042.174p 0.650578mV 560060.545p 0.65798mV 560075.41p 0.695431mV 561003.362p 0.549961mV 561012.949p 0.549829mV 561018.754p 0.576269mV 561065.977p 0.647908mV 562020.168p 0.595276mV 562037.089p 0.618896mV 563023.659p 0.597mV 563042.92p 0.544073mV 563108.995p 0.396605mV 564052.424p 0.656724mV 564069.844p 0.637813mV 566014.832p 0.603614mV 566034.361p 0.654546mV 566038.876p 0.629445mV 566050.869p 0.662924mV 566054.31p 0.662924mV 567016.66p 0.528464mV 567031.785p 0.505313mV 567056.284p 0.482104mV 567059.077p 0.482104mV 567074.892p 0.507635mV 567077.216p 0.532716mV 567134.993p 0.589265mV 567142.389p 0.533839mV 567146.343p 0.558938mV 567167.779p 0.554308mV 567175.404p 0.500063mV 567177.693p 0.500063mV 567220.147p 0.4984mV 568018.682p 0.578715mV 568047.771p 0.638801mV 569000.521p 0.54862mV 569002.043p 0.54862mV 569006.324p 0.575282mV 569044.356p 0.609858mV 569068.127p 0.602056mV 569068.981p 0.602056mV 569070.013p 0.632718mV 570044.651p 0.496474mV 570047.212p 0.468076mV 571001.811p 0.545597mV 571032.888p 0.490447mV 571051.44p 0.431869mV 572003.127p 0.553694mV 572022.806p 0.550496mV 572058.398p 0.469101mV 572072.201p 0.386163mV 573027.678p 0.576003mV 573029.113p 0.576003mV 573044.922p 0.549848mV 573060.472p 0.445831mV 573065.149p 0.419013mV 573077.029p 0.415978mV 573092.576p 0.379468mV 574015.974p 0.474531mV 574023.437p 0.500539mV 574061.681p 0.59588mV 574069.586p 0.568384mV 574072.616p 0.593817mV 574095.063p 0.565658mV 574097.109p 0.565658mV 574103.935p 0.592236mV 574122.26p 0.648487mV 574134.013p 0.653201mV 574138.517p 0.630198mV 574143.198p 0.607929mV 575007.749p 0.526473mV 575009.961p 0.526473mV 575020.84p 0.496409mV 575024.107p 0.496409mV 576037.832p 0.469872mV 576041.201p 0.496218mV 576085.112p 0.508599mV 576102.113p 0.580137mV 576105.782p 0.551408mV 576109.492p 0.551408mV 576116.587p 0.599264mV 576143.622p 0.616498mV 576154.407p 0.614176mV 576190.016p 0.559987mV 576212.935p 0.614283mV 576221.276p 0.616804mV 576234.963p 0.673191mV 576237.152p 0.649702mV 576246.202p 0.657366mV 576250.647p 0.636379mV 576254.278p 0.636379mV 577025.522p 0.63353mV 577034.161p 0.6084mV 577076.894p 0.554625mV 577078.07p 0.554625mV 577096.431p 0.569531mV 577132.058p 0.575645mV 578082.84p 0.688342mV 579014.257p 0.499974mV 579036.208p 0.575232mV 580010.078p 0.54757mV 580015.89p 0.520576mV 580052.45p 0.647258mV 580054.504p 0.647258mV 580079.507p 0.57535mV 580110.013p 0.516324mV 580111.468p 0.516324mV 580138.767p 0.605602mV 580144.444p 0.633831mV 580160.554p 0.645443mV 580166.174p 0.623212mV 580179.4p 0.580676mV 580188.68p 0.642899mV 581016.88p 0.573242mV 581018.382p 0.573242mV 581027.133p 0.574116mV 581034.51p 0.600947mV 581073.931p 0.613422mV 581074.675p 0.613422mV 581077.321p 0.590335mV 581092.133p 0.627742mV 581097.266p 0.606222mV 581101.544p 0.585275mV 582013.764p 0.609465mV 582015.102p 0.63718mV 582023.977p 0.612679mV 582028.242p 0.588772mV 582035.858p 0.59449mV 582057.473p 0.609093mV 582073.963p 0.700186mV 583001.685p 0.553883mV 583002.51p 0.553883mV 583002.566p 0.553883mV 583007.082p 0.526364mV 583020.34p 0.60147mV 583027.235p 0.626635mV 583040.689p 0.652095mV 583045.108p 0.626537mV 583054.606p 0.654255mV 583069.015p 0.688218mV 584006.583p 0.574546mV 584023.95p 0.551684mV 584055.07p 0.588281mV 585019.99p 0.472286mV 585031.047p 0.495mV 585042.692p 0.490466mV 586039.666p 0.406946mV 586047.495p 0.399818mV 587028.175p 0.576312mV 587054.539p 0.54769mV 587056.998p 0.520647mV 587075.833p 0.516286mV 587080.35p 0.488488mV 587082.208p 0.488488mV 587093.266p 0.537227mV 587094.384p 0.537227mV 587130.116p 0.564957mV 587186.711p 0.490868mV 588000.178p 0.548691mV 588007.974p 0.52229mV 589013.604p 0.545731mV 589017.923p 0.571218mV 589042.16p 0.43489mV 590027.645p 0.466156mV 590053.092p 0.477625mV 591037.571p 0.519914mV 591065.792p 0.570932mV 591146.282p 0.453139mV 592028.329p 0.475548mV 592030.897p 0.448812mV 592033.499p 0.448812mV 592046.72p 0.470371mV 592058.019p 0.516257mV 592076.956p 0.498794mV 592080.837p 0.467581mV 593004.431p 0.54976mV 593018.306p 0.578875mV 593030.835p 0.609054mV 594064.002p 0.62883mV 594073.689p 0.689328mV 595017.508p 0.52699mV 595027.921p 0.580849mV 595042.601p 0.503914mV 595068.06p 0.47659mV 595076.811p 0.52509mV 595093.523p 0.490917mV 595102.538p 0.484706mV 595105.554p 0.454821mV 595110.314p 0.476611mV 596004.736p 0.550699mV 596007.346p 0.57822mV 596021.013p 0.555914mV 596040.466p 0.614508mV 596041.172p 0.614508mV 596046.857p 0.590379mV 596060.001p 0.624756mV 596070.579p 0.63151mV 596072.538p 0.63151mV 597002.442p 0.546302mV 597010.925p 0.543591mV 597032.586p 0.591664mV 597121.812p 0.48853mV 598006.032p 0.57855mV 598012.861p 0.551244mV 598019.933p 0.57677mV 598061.364p 0.648637mV 598085.678p 0.681276mV 598089.308p 0.681276mV 598096.151p 0.68948mV 599000.165p 0.547926mV 599017.688p 0.520636mV 599022.044p 0.493841mV 599030.848p 0.492193mV 599031.846p 0.492193mV 599039.18p 0.516973mV 599041.476p 0.541363mV 599051.606p 0.589637mV 599070.149p 0.636127mV 599072.137p 0.636127mV 599078.169p 0.609333mV 599091.081p 0.584204mV 599102.019p 0.639138mV 599106.242p 0.66707mV 600007.198p 0.524165mV 600044.345p 0.493736mV 600046.951p 0.517448mV 600052.417p 0.54077mV 600075.135p 0.54926mV 600101.606p 0.44845mV 601028.594p 0.573827mV 601053.509p 0.604159mV 602007.625p 0.580415mV 602021.992p 0.659689mV 602022.673p 0.659689mV 602035.284p 0.637953mV 603006.18p 0.523211mV 603017.253p 0.577132mV 603033.005p 0.605441mV 603042.728p 0.607578mV 603062.692p 0.668319mV 603071.107p 0.72772mV 604040.314p 0.433051mV 604049.861p 0.4561mV 604063.291p 0.468943mV 605027.009p 0.525954mV 605032.737p 0.551938mV 605042.122p 0.550935mV 605092.732p 0.555083mV 605106.232p 0.534357mV 605107.99p 0.534357mV 606026.433p 0.523367mV 606051.287p 0.65312mV 606058.581p 0.627193mV 606080.235p 0.609747mV 606091.334p 0.562905mV 606100.816p 0.517078mV 606109.333p 0.546434mV 606122.024p 0.5294mV 607028.301p 0.414255mV 608019.819p 0.576513mV 608050.726p 0.659623mV 608054.207p 0.659623mV 608081.247p 0.579024mV 608089.275p 0.557824mV 608117.508p 0.58595mV 608133.417p 0.573524mV 609030.053p 0.497201mV 609044.6p 0.494919mV 610009.851p 0.529124mV 610056.397p 0.535753mV 610057.012p 0.535753mV 610076.832p 0.532716mV 610099.119p 0.527641mV 610104.573p 0.499321mV 610107.718p 0.470874mV 611004.408p 0.551155mV 611021.913p 0.498679mV 612001.87p 0.554354mV 612035.525p 0.638971mV 612049.258p 0.641868mV 612053.922p 0.670263mV 613003.42p 0.547602mV 613015.903p 0.627134mV 613052.826p 0.613865mV 613060.581p 0.621493mV 614001.189p 0.552094mV 614001.3p 0.552094mV 614010.781p 0.60243mV 614042.042p 0.603466mV 614050.615p 0.659938mV 614062.301p 0.71822mV 615010.762p 0.604689mV 615014.024p 0.604689mV 615029.146p 0.579627mV 615058.549p 0.694975mV 615065.276p 0.702496mV 615066.1p 0.702496mV 615068.883p 0.702496mV 616045.476p 0.566124mV 616056.295p 0.51097mV 616056.868p 0.51097mV 616098.174p 0.660399mV 616120.697p 0.593901mV 616131.409p 0.602313mV 616169.524p 0.61303mV 617021.283p 0.550753mV 617021.599p 0.550753mV 617043.578p 0.556023mV 617082.948p 0.621131mV 617091.998p 0.680346mV 617092.826p 0.680346mV 617095.223p 0.710649mV 618011.069p 0.54415mV 618050.073p 0.537372mV 618087.71p 0.496607mV 618090.947p 0.519543mV 619023.72p 0.649787mV 619031.115p 0.650119mV 619032.92p 0.650119mV 619036.916p 0.677383mV 619040.461p 0.705239mV 620001.078p 0.548299mV 620025.217p 0.630819mV 620048.301p 0.58638mV 620052.275p 0.615138mV 621092.222p 0.332656mV 622031.993p 0.501958mV 622091.187p 0.434729mV 623003.523p 0.546262mV 623005.507p 0.571629mV 623032.362p 0.54038mV 623047.623p 0.616259mV 623091.976p 0.544478mV 623110.641p 0.550385mV 623122.2p 0.500478mV 623129.252p 0.475363mV 623167.728p 0.47244mV 623175.669p 0.467653mV 623200.863p 0.473562mV 623201.605p 0.473562mV 624036.94p 0.571214mV 624037.725p 0.571214mV 624094.712p 0.488312mV 624109.108p 0.454656mV 624110.429p 0.42532mV 625019.86p 0.523451mV 626035.259p 0.467667mV 626052.389p 0.438116mV 627002.76p 0.545837mV 627008.121p 0.520181mV 627010.393p 0.547165mV 627029.677p 0.574676mV 627037.733p 0.522656mV 627039.381p 0.522656mV 627075.249p 0.467455mV 627110.133p 0.528234mV 627114.866p 0.528234mV 627115.984p 0.550944mV 627126.237p 0.543853mV 627133.566p 0.514332mV 627135.205p 0.53702mV 627156.516p 0.522171mV 627198.277p 0.53942mV 627213.641p 0.551456mV 627222.837p 0.54199mV 627228.093p 0.511193mV 627239.287p 0.501006mV 628000.088p 0.553881mV 628035.409p 0.628663mV 628044.88p 0.603126mV 629021.421p 0.607368mV 629022.451p 0.607368mV 629041.491p 0.614722mV 629057.643p 0.651389mV 629063.279p 0.682053mV 630004.171p 0.551628mV 630045.614p 0.412765mV 630059.359p 0.404968mV 631018.86p 0.581326mV 631022.347p 0.555778mV 631079.898p 0.361415mV 632003.973p 0.546113mV 632007.687p 0.520603mV 632011.135p 0.547727mV 632025.942p 0.523016mV 632059.729p 0.576612mV 632065.37p 0.6312mV 632094.403p 0.510442mV 632101.189p 0.462519mV 632102.497p 0.462519mV 632125.998p 0.599156mV 632130.304p 0.626232mV 633008.471p 0.573088mV 633054.019p 0.658263mV 634027.089p 0.46649mV 634027.877p 0.46649mV 634055.091p 0.551518mV 634087.288p 0.421283mV 635065.27p 0.647406mV 635078.168p 0.604671mV 636009.357p 0.579797mV 636012.041p 0.605703mV 636014.016p 0.605703mV 636020.535p 0.658249mV 636026.908p 0.632535mV 636054.121p 0.617415mV 637016.942p 0.574693mV 637031.985p 0.65643mV 637033.422p 0.65643mV 637034.582p 0.65643mV 637055.069p 0.591316mV 637085.739p 0.564403mV 637104.689p 0.552905mV 638016.207p 0.574066mV 638024.578p 0.599813mV 639005.963p 0.572945mV 639013.244p 0.598388mV 639017.875p 0.571319mV 639028.029p 0.517908mV 639030.45p 0.491235mV 639038.191p 0.464364mV 639056.134p 0.45782mV 639073.238p 0.421019mV 640035.646p 0.518386mV 640042.856p 0.490325mV 640061.801p 0.374755mV 640066.84p 0.344344mV 641011.354p 0.501503mV 641041.387p 0.495543mV 641042.139p 0.495543mV 641046.213p 0.519172mV 641058.076p 0.565454mV 641081.44p 0.577829mV 641119.688p 0.534316mV 641142.263p 0.490252mV 642017.693p 0.580949mV 642044.115p 0.453238mV 642063.768p 0.555905mV 642108.17p 0.582344mV 642137.366p 0.652592mV 643029.147p 0.467398mV 643046.223p 0.454488mV 643046.436p 0.454488mV 644017.168p 0.579959mV 644030.226p 0.555087mV 644043.99p 0.608657mV 644050.589p 0.5577mV 644057.914p 0.585254mV 644091.032p 0.568494mV 644092.867p 0.568494mV 644096.818p 0.54339mV 644097.686p 0.54339mV 644107.58p 0.546002mV 644114.887p 0.520769mV 644115.638p 0.495508mV 644118.001p 0.495508mV 644167.516p 0.605511mV 644173.366p 0.580595mV 644176.267p 0.608619mV 644183.045p 0.584276mV 644220.617p 0.553187mV 644239.135p 0.535718mV 644241.137p 0.564975mV 644267.302p 0.554298mV 644271.505p 0.583768mV 644281.608p 0.590727mV 645018.199p 0.579209mV 645027.351p 0.581516mV 645052.934p 0.671943mV 645056.83p 0.649894mV 646001.843p 0.55113mV 646003.737p 0.55113mV 646008.61p 0.524307mV 646013.667p 0.550166mV 646036.08p 0.627278mV 646047.04p 0.628423mV 646067.724p 0.690524mV 646071.345p 0.668998mV 647013.898p 0.598601mV 647029.695p 0.571815mV 647038.17p 0.519974mV 648003.448p 0.545708mV 648009.175p 0.572146mV 648029.826p 0.626266mV 648032.869p 0.653555mV 649079.024p 0.576867mV 649089.383p 0.574911mV 649123.397p 0.600244mV 649130.495p 0.655112mV 649134.512p 0.655112mV 649143.696p 0.60677mV 649146.397p 0.635876mV 650002.396p 0.553926mV 650004.877p 0.553926mV 650053.026p 0.512368mV 650059.544p 0.487891mV 650076.169p 0.439498mV 650097.053p 0.434762mV 650110.78p 0.44809mV 651012.416p 0.55186mV 651016.248p 0.524954mV 651044.268p 0.439963mV 651048.115p 0.463462mV 651050.554p 0.486187mV 651055.133p 0.508293mV 651074.57p 0.416551mV 652007.628p 0.580645mV 652008.897p 0.580645mV 652018.544p 0.530441mV 652043.96p 0.455698mV 652071.236p 0.337964mV 653004.3p 0.553618mV 653036.207p 0.633014mV 653056.258p 0.691658mV 653061.32p 0.720904mV 653065.685p 0.698807mV 653065.994p 0.698807mV 654024.815p 0.491823mV 654028.554p 0.464533mV 654058.069p 0.395275mV 655009.499p 0.573938mV 655009.56p 0.573938mV 655047.646p 0.516147mV 655047.878p 0.516147mV 655051.639p 0.542142mV 656009.479p 0.522153mV 656023.823p 0.491585mV 656043.973p 0.429498mV 656046.669p 0.451702mV 657036.183p 0.62672mV 657078.814p 0.64035mV 657081.222p 0.617041mV 657088.003p 0.646603mV 657092.515p 0.676514mV 658020.063p 0.603109mV 658047.622p 0.579028mV 658091.93p 0.678829mV 658099.337p 0.709583mV 659008.142p 0.52675mV 659009.775p 0.52675mV 659016.479p 0.475293mV 659018.71p 0.475293mV 659045.818p 0.521052mV 659052.912p 0.49205mV 659061.066p 0.538016mV 659065.864p 0.560548mV 659074.441p 0.582994mV 659087.464p 0.599166mV 659093.697p 0.570119mV 659094.676p 0.570119mV 659104.812p 0.617587mV 659121.341p 0.717356mV 659124.264p 0.717356mV 660021.626p 0.602272mV 660061.112p 0.552789mV 660084.091p 0.452394mV 660084.769p 0.452394mV 661013.638p 0.551106mV 661054.657p 0.559112mV 661109.01p 0.42685mV 662012.641p 0.494526mV 662016.94p 0.520162mV 662048.04p 0.564857mV 662054.74p 0.537409mV 662068.539p 0.613181mV 662073.266p 0.586056mV 662093.921p 0.638169mV 662129.651p 0.679638mV 663017.937p 0.520249mV 663059.989p 0.447222mV 664033.955p 0.720944mV 664035.319p 0.698514mV 665072.792p 0.625756mV 665075.3p 0.598232mV 665125.98p 0.606193mV 665127.01p 0.606193mV 665249.59p 0.400194mV 666071.564p 0.616804mV 666077.661p 0.645494mV 666093.345p 0.68213mV 667007.836p 0.519379mV 667024.194p 0.438894mV 668001.434p 0.550814mV 668010.798p 0.551038mV 668016.098p 0.524651mV 668029.774p 0.524412mV 668048.731p 0.627331mV 668064.203p 0.601698mV 668073.738p 0.551598mV 668093.931p 0.610956mV 668159.003p 0.581327mV 668163.648p 0.560732mV 668163.696p 0.560732mV 668172.958p 0.571654mV 669003.321p 0.551429mV 669011.023p 0.552361mV 669063.432p 0.444245mV 670019.559p 0.627106mV 670022.863p 0.653327mV 670061.918p 0.569565mV 670077.227p 0.558428mV 671094.874p 0.581035mV 671098.564p 0.551936mV 671113.703p 0.622576mV 671123.055p 0.671086mV 671165.309p 0.60198mV 672014.531p 0.547158mV 672043.27p 0.387157mV 673010.102p 0.604394mV 673014.63p 0.604394mV 673063.601p 0.627999mV 673080.134p 0.595007mV 674014.397p 0.551199mV 674035.785p 0.624764mV 674049.771p 0.677669mV 674067.342p 0.685936mV 675001.26p 0.553644mV 675019.551p 0.531417mV 675062.831p 0.459057mV 675073.372p 0.457496mV 676034.27p 0.556652mV 676094.704p 0.537021mV 676122.567p 0.548561mV 676134.736p 0.551118mV 676153.338p 0.608894mV 676153.635p 0.608894mV 676189.034p 0.605155mV 677034.908p 0.601176mV 677038.813p 0.576336mV 677040.566p 0.55184mV 677070.306p 0.617751mV 677092.248p 0.632773mV 678012.612p 0.552161mV 678017.832p 0.525551mV 678053.676p 0.495292mV 678107.567p 0.536885mV 678159.804p 0.534929mV 679006.065p 0.526267mV 679032.557p 0.558508mV 679038.852p 0.533386mV 679056.949p 0.591052mV 679085.402p 0.709157mV 679089.908p 0.709157mV 679091.494p 0.687142mV 680002.753p 0.553844mV 680039.31p 0.522383mV 680074.395p 0.53964mV 680092.563p 0.530091mV 680130.13p 0.557505mV 680133.974p 0.557505mV 680144.903p 0.601947mV 680163.199p 0.694636mV 680177.792p 0.719163mV 680196.952p 0.676441mV 680202.034p 0.706768mV 681005.081p 0.518382mV 681007.794p 0.518382mV 682004.635p 0.549855mV 682024.902p 0.551246mV 682032.343p 0.551472mV 682041.897p 0.552064mV 682050.407p 0.553032mV 682096.097p 0.58772mV 682110.456p 0.566349mV 682124.94p 0.570935mV 682134.41p 0.576298mV 682155.848p 0.619864mV 682162.686p 0.650756mV 683023.787p 0.493697mV 683027.805p 0.46645mV 683046.866p 0.406093mV 683055.799p 0.398535mV 684040.353p 0.500753mV 684041.515p 0.500753mV 684072.949p 0.440124mV 684085.003p 0.455049mV 685028.315p 0.579473mV 685053.09p 0.504583mV 685118.845p 0.52014mV 685131.386p 0.537284mV 685154.81p 0.575511mV 685166.388p 0.59201mV 685238.433p 0.555215mV 685262.519p 0.570902mV 685262.924p 0.570902mV 685271.249p 0.515008mV 685293.488p 0.401472mV 686007.744p 0.57602mV 686011.195p 0.602146mV 686039.091p 0.63084mV 686053.636p 0.610143mV 686082.819p 0.633058mV 687000.595p 0.552109mV 687037.745p 0.580796mV 687043.379p 0.60737mV 687044.063p 0.60737mV 687049.854p 0.634135mV 687050.456p 0.661252mV 687073.458p 0.617536mV 687075.191p 0.594936mV 687081.697p 0.62492mV 688010.885p 0.603456mV 688053.562p 0.610592mV 688054.162p 0.610592mV 689012.744p 0.601115mV 689025.171p 0.630636mV 690003.044p 0.549972mV 690012.924p 0.600307mV 690094.577p 0.564385mV 690096.908p 0.540668mV 690102.688p 0.517049mV 690116.819p 0.497638mV 690119.087p 0.497638mV 690144.032p 0.475533mV 690146.237p 0.448126mV 690165.738p 0.491206mV 690168.328p 0.491206mV 691042.782p 0.399196mV 691048.785p 0.424073mV 692006.42p 0.527007mV 692101.31p 0.527974mV 692106.817p 0.496574mV 693033.307p 0.705901mV 694009.554p 0.579468mV 694012.743p 0.607103mV 694021.829p 0.610461mV 694028.223p 0.638793mV 694029.83p 0.638793mV 694050.931p 0.734338mV 695000.262p 0.552644mV 695065.743p 0.599907mV 695080.729p 0.687357mV 695084.967p 0.687357mV 696003.026p 0.547526mV 696014.266p 0.546639mV 696079.438p 0.687104mV 696084.498p 0.716891mV 697002.189p 0.548259mV 697019.979p 0.520103mV 697057.848p 0.504611mV 697071.309p 0.46703mV 698000.847p 0.545648mV 698003.512p 0.545648mV 698015.849p 0.62609mV 698045.826p 0.58474mV 698073.809p 0.628267mV 698078.206p 0.659095mV 699003.345p 0.554335mV 699015.548p 0.631793mV 699018.233p 0.631793mV 699025.11p 0.684926mV 699034.831p 0.712398mV 699036.511p 0.688121mV 699046.972p 0.694881mV 700018.08p 0.576267mV 700036.3p 0.633121mV 700048.645p 0.690669mV 700048.88p 0.690669mV 701004.729p 0.553273mV 701058.904p 0.586761mV 701085.416p 0.539314mV 701089.478p 0.539314mV 702006.524p 0.573184mV 702012.198p 0.599215mV 702014.822p 0.599215mV 702028.49p 0.57349mV 702043.438p 0.497612mV 702053.077p 0.499085mV 703010.137p 0.550474mV 703018.013p 0.575377mV 703030.189p 0.597808mV 703031.904p 0.597808mV 703031.933p 0.597808mV 703043.847p 0.543244mV 703069.273p 0.511322mV 703075.639p 0.506563mV 703082.177p 0.477747mV 703087.813p 0.501065mV 704003.077p 0.547642mV 704015.572p 0.57019mV 704019.754p 0.57019mV 704020.364p 0.542474mV 704028.783p 0.567499mV 704030.16p 0.592475mV 704038.98p 0.617567mV 704039.64p 0.617567mV 704058.438p 0.563931mV 704068.653p 0.61813mV 704073.635p 0.592879mV 704097.108p 0.630844mV 704097.588p 0.630844mV 705003.416p 0.550828mV 705006.566p 0.576714mV 705007.1p 0.576714mV 705031.244p 0.495474mV 705032.657p 0.495474mV 705034.77p 0.495474mV 705036.655p 0.520845mV 705047.567p 0.570673mV 705053.714p 0.542866mV 705065.665p 0.512445mV 705066.369p 0.512445mV 705128.632p 0.508181mV 705143.35p 0.484858mV 705148.486p 0.45856mV 705192.335p 0.571797mV 706007.636p 0.524541mV 706026.278p 0.572952mV 706029.002p 0.572952mV 706047.257p 0.568508mV 706069.236p 0.511715mV 706077.323p 0.560838mV 706099.83p 0.552787mV 706161.459p 0.4888mV 707002.121p 0.548622mV 707029.292p 0.519385mV 707066.772p 0.455219mV 708000.626p 0.551972mV 708001.234p 0.551972mV 708001.384p 0.551972mV 708065.313p 0.527246mV 708075.879p 0.576911mV 708077.913p 0.576911mV 708084.779p 0.601682mV 708097.77p 0.5724mV 708101.519p 0.598503mV 708112.382p 0.651298mV 709024.453p 0.605527mV 709035.508p 0.636996mV 709037.545p 0.636996mV 709065.802p 0.607913mV 709068.441p 0.607913mV 710005.247p 0.571963mV 710015.426p 0.569619mV 710029.305p 0.568131mV 710037.041p 0.567454mV 710069.942p 0.570102mV 710077.099p 0.519957mV 710121.4p 0.55242mV 710145.91p 0.47773mV 710151.127p 0.45194mV 710164.133p 0.451508mV 710165.309p 0.476857mV 710185.777p 0.468003mV 711014.986p 0.604078mV 711035.296p 0.478256mV 711046.153p 0.479592mV 711046.926p 0.479592mV 711047.143p 0.479592mV 711050.246p 0.453419mV 712069.428p 0.596741mV 712099.825p 0.582578mV 712119.015p 0.632069mV 712120.026p 0.605502mV 712127.142p 0.579453mV 712134.535p 0.606427mV 712189.838p 0.491575mV 712196.799p 0.545425mV 712212.003p 0.519462mV 712216.66p 0.492751mV 712222.674p 0.465852mV 712232.717p 0.463501mV 712233.475p 0.463501mV 712254.404p 0.558451mV 712278.77p 0.411108mV 713000.128p 0.552487mV 713037.957p 0.423925mV 714013.826p 0.547069mV 714043.466p 0.547318mV 714095.582p 0.402081mV 715009.841p 0.521153mV 716013.763p 0.494328mV 716048.054p 0.406338mV 716062.673p 0.420244mV 717005.976p 0.522766mV 717009.694p 0.522766mV 717025.049p 0.627007mV 717026.424p 0.627007mV 717049.667p 0.631114mV 718036.409p 0.425157mV 719058.032p 0.546768mV 719065.52p 0.551416mV 719070.555p 0.527303mV 719120.044p 0.608735mV 720006.097p 0.524109mV 720010.33p 0.550118mV 720064.438p 0.653153mV 720066.936p 0.628727mV 720090.913p 0.620542mV 720091.353p 0.620542mV 721030.182p 0.611838mV 722021.034p 0.49394mV 722034.262p 0.440507mV 722034.789p 0.440507mV 722043.166p 0.437652mV 723008.685p 0.581188mV 723012.974p 0.608421mV 724037.566p 0.637118mV 724053.812p 0.618011mV 724053.875p 0.618011mV 725014.986p 0.548439mV 725068.538p 0.551064mV 725096.394p 0.533135mV 726043.387p 0.43912mV 727047.969p 0.581132mV 727059.797p 0.635643mV 727070.602p 0.720359mV 727074.441p 0.720359mV 728003.608p 0.549032mV 728007.853p 0.52158mV 728016.547p 0.571747mV 728096.542p 0.570283mV 728142.029p 0.514272mV 728189.009p 0.508362mV 728197.931p 0.510775mV 728212.325p 0.486537mV 728217.625p 0.512649mV 729003.669p 0.552522mV 729006.158p 0.578443mV 729007.466p 0.578443mV 729012.276p 0.551704mV 729049.956p 0.520472mV 729070.742p 0.590499mV 729094.07p 0.693662mV 729098.042p 0.720878mV 729099.917p 0.720878mV 729108.394p 0.725561mV 729112.089p 0.703587mV 730008.811p 0.579528mV 730010.978p 0.607259mV 730021.196p 0.663398mV 730029.984p 0.639665mV 730116.448p 0.441256mV 730125.422p 0.442451mV 731004.577p 0.547604mV 731020.727p 0.496421mV 731035.325p 0.574896mV 731036.243p 0.574896mV 731039.973p 0.574896mV 731040.586p 0.600819mV 731074.205p 0.606074mV 732032.005p 0.493134mV 732036.605p 0.517607mV 733020.018p 0.599875mV 733032.96p 0.60037mV 733069.328p 0.585516mV 733094.721p 0.632321mV 734005.386p 0.578164mV 734007.705p 0.578164mV 734024.005p 0.608511mV 734043.753p 0.566254mV 734045.475p 0.543141mV 734056.737p 0.549412mV 734082.074p 0.644237mV 735000.075p 0.552237mV 735000.178p 0.552237mV 735019.666p 0.581493mV 735042.475p 0.510662mV 735050.746p 0.460921mV 735057.233p 0.435497mV 735062.722p 0.4095mV 737027.04p 0.571376mV 737037.482p 0.622937mV 737061.14p 0.600983mV 737062.986p 0.600983mV 737075.933p 0.688024mV 737080.841p 0.665888mV 737085.01p 0.644757mV 738012.394p 0.603829mV 738012.514p 0.603829mV 738041.565p 0.56326mV 738076.931p 0.611876mV 738084.799p 0.641349mV 739004.114p 0.552555mV 739031.759p 0.557931mV 739073.094p 0.568164mV 739084.874p 0.572794mV 739101.29p 0.529961mV 739155.465p 0.510434mV 739191.302p 0.514758mV 740001.35p 0.551612mV 740048.012p 0.578295mV 740058.162p 0.527885mV 741022.093p 0.490223mV 741051.703p 0.474219mV 741060.224p 0.464332mV 742000.604p 0.545894mV 742015.4p 0.521483mV 742022.666p 0.495861mV 742074.361p 0.485621mV 742084.528p 0.425612mV 742088.367p 0.39498mV 743005.37p 0.519301mV 743014.117p 0.492328mV 743020.088p 0.542943mV 743062.104p 0.581487mV 743105.511p 0.596177mV 743116.735p 0.542689mV 743125.14p 0.542364mV 743125.555p 0.542364mV 743126.621p 0.542364mV 743132.697p 0.515627mV 743136.624p 0.541519mV 743192.42p 0.684948mV 743194.686p 0.684948mV 744043.901p 0.495455mV 744045.5p 0.520128mV 744081.481p 0.419213mV 745018.365p 0.580862mV 745028.748p 0.58468mV 745030.014p 0.560813mV 745034.505p 0.560813mV 745041.29p 0.513635mV 745064.878p 0.469468mV 745079.474p 0.44473mV 745087.775p 0.495561mV 746028.252p 0.530118mV 746062.002p 0.504567mV 746088.511p 0.473289mV 746106.22p 0.569191mV 746130.172p 0.476456mV 746147.9p 0.438566mV 747004.324p 0.549803mV 747010.933p 0.601197mV 747015.527p 0.574383mV 747052.487p 0.49269mV 747087.625p 0.501552mV 748014.317p 0.548213mV 748047.114p 0.464825mV 748080.935p 0.468917mV 748083.719p 0.468917mV 748084.933p 0.468917mV 748086.475p 0.489766mV 748089.648p 0.489766mV 749000.823p 0.55406mV 749005.031p 0.52669mV 749020.266p 0.444076mV 749038.444p 0.409855mV 750018.511p 0.472973mV 750052.663p 0.594381mV 750066.104p 0.566115mV 750070.59p 0.592246mV 750107.834p 0.567934mV 750116.588p 0.56927mV 750131.11p 0.545518mV 750155.21p 0.578378mV 750161.728p 0.606167mV 751027.23p 0.576371mV 751034.307p 0.603766mV 751036.115p 0.578694mV 751065.567p 0.538608mV 751086.763p 0.600734mV 752008.743p 0.573279mV 752010.752p 0.598447mV 752032.053p 0.648605mV 752048.851p 0.677163mV 753013.778p 0.606962mV 753020.868p 0.555084mV 753037.527p 0.531349mV 753096.44p 0.417494mV 754065.94p 0.525087mV 754081.412p 0.547807mV 754112.098p 0.484691mV 754117.479p 0.508914mV 755064.24p 0.476505mV 756002.758p 0.551154mV 756023.173p 0.500061mV 756039.492p 0.420475mV 757000.016p 0.54652mV 757006.805p 0.519626mV 757031.48p 0.434555mV 757033.026p 0.434555mV 758011.497p 0.55237mV 758025.772p 0.475967mV 759018.089p 0.570348mV 759021.042p 0.595594mV 759046.222p 0.566043mV 759054.535p 0.591828mV 759068.106p 0.670452mV 759072.595p 0.697607mV 760037.435p 0.512693mV 760072.159p 0.570158mV 760095.982p 0.633495mV 760096.166p 0.633495mV 760105.096p 0.629149mV 760112.954p 0.601615mV 760113.765p 0.601615mV 760135.03p 0.62623mV 761002.615p 0.547597mV 761063.345p 0.37677mV 762073.513p 0.425506mV 763024.864p 0.551385mV 763027.236p 0.524837mV 763043.887p 0.497254mV 763051.168p 0.494585mV 763055.634p 0.519193mV 763067.943p 0.514951mV 763091.418p 0.526688mV 763115.442p 0.637673mV 763146.438p 0.627338mV 763167.721p 0.632147mV 763168.585p 0.632147mV 763182.861p 0.615879mV 763192.808p 0.676998mV 763193.549p 0.676998mV 764006.455p 0.573654mV 764008.717p 0.573654mV 764010.828p 0.59881mV 764011.463p 0.59881mV 764026.416p 0.622873mV 764045.215p 0.677895mV 764053.197p 0.654215mV 764053.463p 0.654215mV 764054.87p 0.654215mV 765000.721p 0.55265mV 765014.566p 0.602452mV 765023.589p 0.600332mV 765044.677p 0.706614mV 765045.665p 0.682169mV 765073.576p 0.676509mV 766009.16p 0.524803mV 766028.186p 0.571719mV 766048.992p 0.618329mV 767005.434p 0.580807mV 767034.082p 0.609961mV 767050.169p 0.614653mV 767053.075p 0.614653mV 767061.219p 0.618399mV 767061.508p 0.618399mV 767069.014p 0.594833mV 767089.901p 0.660701mV 767093.072p 0.638998mV 767096.556p 0.618109mV 768000.902p 0.549277mV 768010.082p 0.547517mV 768023.376p 0.545385mV 768023.495p 0.545385mV 768029.227p 0.570434mV 768050.697p 0.538529mV 768068.237p 0.509973mV 768068.395p 0.509973mV 768072.776p 0.482855mV 768079.627p 0.508137mV 768087.223p 0.504935mV 768108.788p 0.547662mV 768124.652p 0.514002mV 768133.17p 0.560144mV 768139.021p 0.582998mV 768144.453p 0.605925mV 768163.473p 0.649012mV 768183.776p 0.701852mV 769009.806p 0.573944mV 769010.345p 0.599316mV 769043.129p 0.597779mV 769058.815p 0.520077mV 769067.307p 0.521087mV 769101.459p 0.493226mV 769121.477p 0.433579mV 769129.237p 0.456206mV 770007.916p 0.573577mV 770009.543p 0.573577mV 770024.332p 0.54527mV 770031.375p 0.596266mV 770071.921p 0.6532mV 770076.994p 0.682284mV 771004.318p 0.552957mV 771016.17p 0.634145mV 771020.655p 0.661677mV 771025.975p 0.637133mV 771028.477p 0.637133mV 771045.786p 0.65067mV 772036.385p 0.522959mV 772036.873p 0.522959mV 772048.712p 0.520655mV 772060.108p 0.488884mV 772067.447p 0.512441mV 772110.943p 0.505639mV 772113.47p 0.505639mV 773029.822p 0.473788mV 773045.451p 0.523787mV 773059.797p 0.520861mV 773061.198p 0.5456mV 773119.955p 0.497667mV 773133.454p 0.460166mV 774007.33p 0.521386mV 774013.818p 0.548761mV 774018.297p 0.575963mV 774032.231p 0.605536mV 774042.668p 0.556392mV 774073.69p 0.461351mV 774098.321p 0.377082mV 775017.685p 0.572542mV 775032.335p 0.545711mV 775074.454p 0.651664mV 775080.731p 0.654534mV 775083.163p 0.654534mV 775112.06p 0.572269mV 775112.229p 0.572269mV 775119.255p 0.550616mV 776003.076p 0.546892mV 776006.361p 0.574584mV 776015.684p 0.577462mV 776016.24p 0.577462mV 776017.442p 0.577462mV 776018.011p 0.577462mV 776020.972p 0.552682mV 776021.704p 0.552682mV 776057.2p 0.589431mV 776093.348p 0.62842mV 777012.469p 0.601749mV 777079.119p 0.4907mV 777085.43p 0.439672mV 777104.019p 0.411414mV 777112.741p 0.353875mV 778079.262p 0.589596mV 778081.904p 0.565973mV 778096.642p 0.60119mV 778111.506p 0.639505mV 778113.617p 0.639505mV 779031.416p 0.66628mV 779049.776p 0.701472mV 780003.691p 0.554292mV 780010.178p 0.554371mV 780017.271p 0.527944mV 780024.093p 0.501544mV 780060.941p 0.492553mV 780093.857p 0.525545mV 781014.253p 0.602926mV 781021.327p 0.606291mV 782022.049p 0.545159mV 782034.208p 0.491831mV 782053.471p 0.434207mV 782064.26p 0.480453mV 782078.409p 0.493417mV 783019.398p 0.581004mV 783029.001p 0.530438mV 783048.223p 0.482096mV 784016.084p 0.522206mV 784044.571p 0.485533mV 786008.307p 0.578105mV 786032.263p 0.506336mV 786041.304p 0.561299mV 786057.331p 0.643425mV 786065.042p 0.699837mV 786081.743p 0.685328mV 787022.641p 0.605304mV 787038.65p 0.583654mV 787065.592p 0.653204mV 788021.427p 0.550675mV 788025.278p 0.576875mV 788067.228p 0.634542mV 788071.355p 0.663326mV 788084.184p 0.722408mV 789013.41p 0.550778mV 789017.815p 0.578191mV 789018.834p 0.578191mV 789032.047p 0.502921mV 789050.477p 0.506115mV 789061.184p 0.453168mV 789064.548p 0.453168mV 789069.213p 0.478789mV 789091.787p 0.546967mV 789118.994p 0.559007mV 789122.371p 0.53046mV 789129.678p 0.554458mV 789143.28p 0.573829mV 789144.691p 0.573829mV 789151.01p 0.569636mV 789166.906p 0.643908mV 789195.385p 0.702265mV 789195.501p 0.702265mV 789202.889p 0.679975mV 790030.498p 0.538327mV 790056.134p 0.451853mV 791021.806p 0.547732mV 791043.29p 0.548227mV 791044.569p 0.548227mV 791064.546p 0.443502mV 791072.283p 0.441442mV 791077.638p 0.413004mV 791082.005p 0.436337mV 792002.37p 0.551527mV 792042.731p 0.555112mV 792057.556p 0.529185mV 792061.837p 0.502939mV 792064.024p 0.502939mV 792089.625p 0.473144mV 792096.11p 0.522142mV 792100.961p 0.49355mV 792114.006p 0.54055mV 792136.186p 0.49758mV 794066.485p 0.691974mV 794066.775p 0.691974mV 794070.3p 0.720608mV 794084.449p 0.780271mV 795002.2p 0.552681mV 795002.939p 0.552681mV 795007.846p 0.525809mV 795009.724p 0.525809mV 795025.205p 0.469836mV 796060.57p 0.517355mV 796066.624p 0.492303mV 796081.161p 0.520864mV 796098.252p 0.54793mV 796100.178p 0.521359mV 796101.847p 0.521359mV 796125.812p 0.544308mV 796138.033p 0.48929mV 796183.652p 0.606134mV 796235.911p 0.524886mV 796242.305p 0.550579mV 796297.722p 0.620342mV 796297.768p 0.620342mV 796306.051p 0.619092mV 796317.486p 0.567262mV 796344.625p 0.706065mV 796354.347p 0.713401mV 797008.833p 0.57654mV 797014.318p 0.601448mV 797041.632p 0.548121mV 797055.418p 0.525071mV 797057.017p 0.525071mV 797067.525p 0.473523mV 797110.532p 0.544039mV 797139.466p 0.506059mV 797142.32p 0.529278mV 797143.777p 0.529278mV 797174.34p 0.615095mV 797182.273p 0.662959mV 797192.94p 0.71321mV 797197.917p 0.739579mV 797206.084p 0.690264mV 797220.065p 0.676437mV 797222.793p 0.676437mV 798000.744p 0.551665mV 798005.226p 0.526751mV 798038.778p 0.478487mV 798050.682p 0.450001mV 798054.478p 0.450001mV 798063.437p 0.445325mV 798075.612p 0.512268mV 798087.579p 0.450856mV 798089.458p 0.450856mV 799000.472p 0.550794mV 799005.457p 0.577099mV 799059.381p 0.477681mV 799109.393p 0.464351mV 800007.752p 0.581201mV 800014.616p 0.608936mV 800038.515p 0.540433mV 800056.243p 0.549582mV 800085.961p 0.506821mV 800133.754p 0.467604mV 801017.29p 0.579596mV 801038.266p 0.584969mV 801043.155p 0.613171mV 801050.914p 0.670327mV 802077.721p 0.497614mV 803002.763p 0.546796mV 803052.4p 0.442311mV 804027.071p 0.572615mV 804027.197p 0.572615mV 805000.318p 0.549971mV 806057.698p 0.625135mV 806089.276p 0.742309mV 807001.775p 0.554355mV 807008.473p 0.57997mV 807022.171p 0.657642mV 807057.96p 0.595851mV 807065.333p 0.605728mV 808011.173p 0.547789mV 808020.028p 0.548296mV 808038.511p 0.521961mV 808049.21p 0.574206mV 808049.737p 0.574206mV 808063.408p 0.547204mV 808095.539p 0.624738mV 808099.909p 0.624738mV 808110.605p 0.706192mV 808122.834p 0.711457mV 808124.414p 0.711457mV 808130.327p 0.668497mV 809012.721p 0.543726mV 809027.324p 0.56678mV 809124.068p 0.609681mV 809124.42p 0.609681mV 809188.942p 0.496952mV 809190.46p 0.46751mV 810057.64p 0.576515mV 810069.819p 0.630357mV 811008.433p 0.526508mV 811025.51p 0.52104mV 811055.322p 0.614283mV 811089.147p 0.669337mV 812069.666p 0.613726mV 812081.92p 0.534394mV 812085.578p 0.560985mV 812105.474p 0.614365mV 812116.324p 0.615633mV 812130.256p 0.593657mV 813010.228p 0.551048mV 813032.601p 0.496289mV 813067.116p 0.618739mV 813077.152p 0.616611mV 813084.609p 0.58968mV 813091.935p 0.589572mV 813112.867p 0.48704mV 813133.326p 0.433405mV 814006.267p 0.522576mV 815068.627p 0.550835mV 815094.381p 0.557181mV 816033.041p 0.551295mV 816040.175p 0.552532mV 816042.503p 0.552532mV 816061.862p 0.502521mV 816092.259p 0.390912mV 817009.494p 0.525819mV 817021.168p 0.494843mV 817071.875p 0.576331mV 817105.292p 0.648493mV 817109.566p 0.648493mV 817111.764p 0.622241mV 817118.554p 0.596618mV 817168.311p 0.563124mV 817204.605p 0.552722mV 817242.056p 0.574829mV 817249.479p 0.552833mV 817254.212p 0.583036mV 817264.346p 0.539679mV 818022.732p 0.448957mV 818046.174p 0.36116mV 819009.682p 0.523012mV 819057.325p 0.558018mV 819065.544p 0.500462mV 819070.271p 0.471592mV 820001.636p 0.552854mV 820032.895p 0.496242mV 820059.86p 0.510089mV 821044.089p 0.442081mV 821068.039p 0.347549mV 822009.148p 0.576079mV 822011.692p 0.602295mV 822020.926p 0.655383mV 822044.062p 0.60957mV 822044.976p 0.60957mV 822052.815p 0.61577mV 822068.383p 0.706559mV 823007.21p 0.578579mV 823023.694p 0.658265mV 823027.946p 0.632964mV 823034.309p 0.60838mV 823037.465p 0.636855mV 823057.057p 0.650055mV 824020.587p 0.554578mV 824036.585p 0.532896mV 824038.792p 0.532896mV 824075.407p 0.656506mV 824086.409p 0.665532mV 825022.828p 0.495632mV 825041.825p 0.544385mV 825053.313p 0.593729mV 825059.489p 0.565914mV 825080.23p 0.532984mV 825093.867p 0.529259mV 825122.952p 0.569689mV 825163.762p 0.667616mV 825164.117p 0.667616mV 825169.06p 0.64301mV 825172.958p 0.619202mV 825178.573p 0.596041mV 825181.382p 0.625604mV 825190.475p 0.581443mV 825198.029p 0.611932mV 825208.798p 0.569998mV 826025.812p 0.524402mV 826049.711p 0.528554mV 827003.691p 0.549276mV 827046.742p 0.471455mV 827061.634p 0.493413mV 827113.988p 0.466036mV 828012.431p 0.596888mV 828016.245p 0.569925mV 828040.401p 0.596498mV 828054.271p 0.59803mV 828056.401p 0.573095mV 828063.893p 0.548481mV 828089.917p 0.477383mV 828097.148p 0.531365mV 828121.141p 0.611596mV 828129.684p 0.58616mV 828150.894p 0.570158mV 828163.326p 0.576625mV 828177.173p 0.612932mV 828180.884p 0.590522mV 828196.724p 0.629623mV 829008.902p 0.572843mV 829011.467p 0.547285mV 829061.042p 0.499905mV 829075.145p 0.579405mV 829076.929p 0.579405mV 830038.609p 0.519186mV 830055.056p 0.566107mV 830056.989p 0.566107mV 830082.821p 0.478998mV 831024.885p 0.444583mV 832021.999p 0.599289mV 832042.772p 0.544226mV 832086.016p 0.52524mV 832100.455p 0.609686mV 832102.44p 0.609686mV 832119.83p 0.642931mV 832128.42p 0.649607mV 832129.913p 0.649607mV 832133.83p 0.679937mV 832139.626p 0.659009mV 833032.64p 0.665586mV 834046.636p 0.522823mV 834068.584p 0.464165mV 834078.272p 0.458012mV 835009.621p 0.578631mV 835032.696p 0.558063mV 835048.526p 0.590657mV 835057.296p 0.595204mV 835060.308p 0.62422mV 835064.832p 0.62422mV 835069.875p 0.653481mV 835089.92p 0.61897mV 836013.962p 0.549261mV 836017.105p 0.523592mV 836020.888p 0.550585mV 836051.024p 0.445975mV 836054.253p 0.445975mV 836057.498p 0.41871mV 836064.004p 0.443417mV 836067.718p 0.414774mV 836069.914p 0.414774mV 837020.287p 0.55231mV 837025.118p 0.578203mV 837027.265p 0.578203mV 837033.913p 0.551435mV 837049.83p 0.47152mV 837054.341p 0.497127mV 839039.979p 0.371503mV 840007.156p 0.579109mV 840061.21p 0.505049mV 840095.081p 0.457755mV 841010.945p 0.600629mV 841034.386p 0.658077mV 841043.127p 0.716135mV 842024.927p 0.502779mV 842040.079p 0.449125mV 842043.362p 0.449125mV 842052.653p 0.49861mV 842064.489p 0.493566mV 842067.281p 0.464244mV 843084.039p 0.542611mV 843096.036p 0.531335mV 843100.879p 0.562176mV 843107.298p 0.592923mV 843110.02p 0.623727mV 844043.47p 0.553955mV 844086.237p 0.655855mV 844086.567p 0.655855mV 845004.931p 0.554247mV 845007.278p 0.529214mV 845032.56p 0.562517mV 845037.69p 0.590834mV 845044.131p 0.619222mV 845059.909p 0.601764mV 845094.735p 0.553976mV 846014.603p 0.551985mV 846016.94p 0.578037mV 846017.166p 0.578037mV 846033.51p 0.498553mV 846046.103p 0.470326mV 846081.213p 0.530817mV 846115.068p 0.581727mV 846129.687p 0.625542mV 846132.022p 0.595782mV 846138.719p 0.566423mV 846143.703p 0.537315mV 846179.071p 0.59624mV 846200.353p 0.615933mV 846228.374p 0.643711mV 846240.792p 0.676259mV 846253.51p 0.683739mV 847010.556p 0.552542mV 847011.026p 0.552542mV 847026.474p 0.631425mV 847032.865p 0.658188mV 847037.822p 0.685446mV 848020.458p 0.496189mV 848021.913p 0.496189mV 848028.687p 0.521566mV 848064.492p 0.425047mV 849041.798p 0.604965mV 849059.701p 0.587256mV 850000.792p 0.552322mV 850008.584p 0.578185mV 850028.661p 0.630415mV 850052.725p 0.666566mV 851001.303p 0.550476mV 851017.543p 0.52809mV 851022.38p 0.50323mV 851046.785p 0.481857mV 851077.133p 0.533824mV 851115.952p 0.527602mV 851123.37p 0.553129mV 851158.652p 0.516906mV 851168.258p 0.459973mV 851190.896p 0.466433mV 852010.413p 0.552468mV 852013.094p 0.552468mV 852016.311p 0.526262mV 852027.088p 0.526413mV 852028.123p 0.526413mV 852062.527p 0.607927mV 852171.638p 0.491297mV 852203.324p 0.474104mV 852215.658p 0.434386mV 852219.003p 0.434386mV 853000.745p 0.548079mV 853001.347p 0.548079mV 853001.616p 0.548079mV 853008.32p 0.521403mV 853041.761p 0.382767mV 854022.845p 0.655128mV 854026.359p 0.630668mV 854043.43p 0.71825mV 855020.828p 0.551139mV 855031.823p 0.606342mV 855032.249p 0.606342mV 855038.76p 0.581516mV 855039.836p 0.581516mV 855059.258p 0.537969mV 855060.464p 0.566872mV 855086.235p 0.555375mV 855107.42p 0.621805mV 855116.547p 0.630631mV 855119.586p 0.630631mV 856000.371p 0.550386mV 856002.343p 0.550386mV 856007.546p 0.575548mV 856040.644p 0.546782mV 856058.269p 0.521359mV 856065.606p 0.574182mV 856075.0p 0.574267mV 856092.403p 0.655202mV 856095.482p 0.630293mV 856099.419p 0.630293mV 856132.21p 0.574969mV 856134.035p 0.574969mV 856137.897p 0.553477mV 856147.31p 0.510882mV 856194.606p 0.570376mV 856220.949p 0.537655mV 856221.583p 0.537655mV 856240.306p 0.500686mV 856242.652p 0.500686mV 856250.747p 0.559875mV 856253.702p 0.559875mV 856267.494p 0.4911mV 856269.555p 0.4911mV 856275.241p 0.49668mV 856284.389p 0.472495mV 856306.176p 0.397711mV 856308.293p 0.397711mV 857012.841p 0.598215mV 857021.224p 0.59712mV 857039.481p 0.676395mV 858000.033p 0.548272mV 858005.189p 0.574646mV 858022.729p 0.549008mV 858067.098p 0.634957mV 858079.62p 0.586425mV 858100.266p 0.627977mV 858115.068p 0.616075mV 859049.189p 0.567025mV 859056.174p 0.565683mV 859059.396p 0.565683mV 859064.813p 0.591335mV 859074.534p 0.590427mV 859086.455p 0.618009mV 859103.81p 0.64981mV 860028.361p 0.572454mV 860032.937p 0.546123mV 860036.683p 0.519934mV 860047.468p 0.467317mV 861012.578p 0.548933mV 861027.454p 0.522533mV 861039.964p 0.522074mV 861068.653p 0.462499mV 861078.735p 0.456815mV 861089.15p 0.501279mV 861103.648p 0.461002mV 862047.785p 0.743782mV 863007.691p 0.520897mV 863019.487p 0.522003mV 863043.69p 0.495511mV 863046.963p 0.46843mV 865030.658p 0.557094mV 865062.587p 0.508159mV 865089.348p 0.535766mV 865104.002p 0.507585mV 865106.139p 0.480558mV 865147.286p 0.512794mV 866013.637p 0.553851mV 867007.571p 0.526064mV 867013.734p 0.552627mV 867017.063p 0.579039mV 867017.289p 0.579039mV 867030.864p 0.606355mV 867052.719p 0.559518mV 867057.838p 0.535539mV 867083.63p 0.571455mV 867089.941p 0.59911mV 867107.025p 0.554063mV 867150.211p 0.548102mV 867185.008p 0.588076mV 867199.25p 0.644067mV 868028.689p 0.575799mV 868056.192p 0.629803mV 869023.527p 0.556142mV 869033.607p 0.558078mV 869052.352p 0.616462mV 869058.965p 0.59231mV 869097.517p 0.45442mV 869119.016p 0.507189mV 869122.194p 0.47966mV 869129.631p 0.451878mV 869145.93p 0.387298mV 870054.374p 0.553826mV 870096.758p 0.574841mV 870115.138p 0.576754mV 870119.397p 0.576754mV 870124.957p 0.551564mV 870148.36p 0.532605mV 871032.61p 0.595088mV 871057.272p 0.566645mV 871062.672p 0.592393mV 871113.858p 0.663732mV 872011.698p 0.601215mV 872012.421p 0.601215mV 872039.907p 0.627787mV 872050.829p 0.554882mV 872063.894p 0.559976mV 872134.245p 0.596989mV 872143.164p 0.551618mV 872177.532p 0.442482mV 872232.502p 0.499919mV 873063.463p 0.595721mV 873090.099p 0.601533mV 873130.533p 0.57508mV 873144.57p 0.635999mV 873145.313p 0.666788mV 873146.306p 0.666788mV 874027.544p 0.463338mV 874045.466p 0.558873mV 874046.723p 0.558873mV 874051.994p 0.582096mV 874066.976p 0.547899mV 874080.832p 0.514896mV 874100.159p 0.502994mV 874114.562p 0.494635mV 875011.306p 0.600366mV 875013.571p 0.600366mV 875066.714p 0.649667mV 876004.564p 0.551492mV 876036.84p 0.464791mV 876050.364p 0.428704mV 877020.188p 0.554608mV 877029.921p 0.52959mV 877032.425p 0.504602mV 877059.698p 0.481761mV 877063.099p 0.507588mV 877088.262p 0.527135mV 877100.491p 0.495204mV 877136.596p 0.49888mV 877156.167p 0.530558mV 878011.021p 0.597854mV 878014.718p 0.597854mV 878017.893p 0.570897mV 878048.276p 0.568573mV 878075.002p 0.510265mV 878075.359p 0.510265mV 878102.087p 0.579912mV 878121.362p 0.573786mV 878127.434p 0.599518mV 878162.224p 0.517994mV 878174.388p 0.514882mV 878205.808p 0.468306mV 879001.216p 0.547312mV 879015.43p 0.569735mV 879017.166p 0.569735mV 879018.847p 0.569735mV 879029.639p 0.568048mV 879036.065p 0.619162mV 879042.737p 0.645059mV 879050.441p 0.64565mV 879074.055p 0.654374mV 880010.928p 0.606359mV 880023.496p 0.60788mV 880025.837p 0.635332mV 880042.44p 0.667823mV 881028.473p 0.518287mV 881029.419p 0.518287mV 881039.147p 0.51548mV 881049.55p 0.564053mV 881073.584p 0.528089mV 882001.714p 0.545625mV 882022.896p 0.593224mV 882033.882p 0.538312mV 882055.066p 0.56064mV 882088.159p 0.615263mV 882102.433p 0.647648mV 883011.8p 0.554148mV 883046.797p 0.587674mV 883104.869p 0.629024mV 883116.509p 0.610198mV 883126.432p 0.617385mV 884042.382p 0.544174mV 884067.766p 0.567222mV 884076.133p 0.512697mV 884078.156p 0.512697mV 884080.926p 0.485426mV 884081.465p 0.485426mV 884085.407p 0.510562mV 884094.227p 0.48268mV 885034.472p 0.601388mV 885041.272p 0.603621mV 885048.989p 0.579105mV 885053.591p 0.554952mV 885069.566p 0.588316mV 885090.191p 0.629587mV 885092.439p 0.629587mV 885100.661p 0.63804mV 885101.506p 0.63804mV 885103.77p 0.63804mV 886011.128p 0.54714mV 886035.544p 0.571395mV 886048.151p 0.624676mV 886053.683p 0.599012mV 886060.719p 0.548983mV 886079.264p 0.474718mV 886091.289p 0.50312mV 886099.683p 0.476985mV 886103.818p 0.450555mV 887007.588p 0.577841mV 887016.023p 0.576568mV 887036.283p 0.628717mV 887051.378p 0.659595mV 887052.761p 0.659595mV 888000.341p 0.547546mV 888006.911p 0.572723mV 888026.652p 0.674915mV 888028.4p 0.674915mV 889021.521p 0.604282mV 889060.333p 0.51458mV 889081.769p 0.577428mV 889091.772p 0.530457mV 889109.958p 0.564666mV 889130.035p 0.602432mV 889158.189p 0.592015mV 889159.699p 0.592015mV 889167.91p 0.601086mV 889213.483p 0.568871mV 889225.874p 0.608913mV 889228.982p 0.608913mV 890063.066p 0.571874mV 890093.174p 0.59155mV 890122.877p 0.461272mV 890124.238p 0.461272mV 890125.714p 0.490967mV 890174.958p 0.421646mV 890176.735p 0.445423mV 890177.627p 0.445423mV 891024.757p 0.55638mV 891050.019p 0.509611mV 891076.521p 0.591193mV 891082.014p 0.565035mV 891085.221p 0.53914mV 891088.29p 0.53914mV 891099.448p 0.487473mV 891100.517p 0.46137mV 891110.671p 0.513173mV 891178.63p 0.543569mV 891201.476p 0.542311mV 892022.325p 0.597493mV 892049.429p 0.51844mV 892062.887p 0.54303mV 892085.266p 0.62049mV 892090.717p 0.647678mV 892092.472p 0.647678mV 893017.983p 0.522102mV 893038.759p 0.57472mV 893072.513p 0.551263mV 893096.906p 0.534346mV 893099.0p 0.534346mV 893114.289p 0.567543mV 893150.185p 0.646087mV 894009.354p 0.520495mV 894018.339p 0.519612mV 894022.663p 0.545051mV 894040.998p 0.592802mV 894041.646p 0.592802mV 894044.571p 0.592802mV 894054.0p 0.643218mV 894084.98p 0.70268mV 895016.531p 0.471251mV 895026.757p 0.416935mV 895030.057p 0.441488mV 896006.804p 0.526987mV 896015.706p 0.527228mV 896025.292p 0.52656mV 897007.563p 0.51862mV 897017.165p 0.463973mV 897026.801p 0.513068mV 897057.278p 0.440413mV 897060.561p 0.40943mV 898001.903p 0.547977mV 898009.29p 0.57456mV 898049.11p 0.5235mV 898076.68p 0.468458mV 898086.641p 0.412722mV 898093.367p 0.436445mV 899018.377p 0.573752mV 899047.193p 0.472131mV 899068.903p 0.417233mV 899077.228p 0.465145mV 900005.765p 0.525223mV 900005.818p 0.525223mV 900019.474p 0.523287mV 901012.53p 0.498474mV 901014.777p 0.498474mV 901047.155p 0.358538mV 902007.431p 0.521728mV 902014.695p 0.549166mV 902018.395p 0.523782mV 902024.912p 0.498393mV 902037.259p 0.473551mV 902055.794p 0.417278mV 902062.903p 0.440885mV 902073.067p 0.433422mV 903013.248p 0.599558mV 903036.621p 0.627045mV 903056.578p 0.583975mV 903056.914p 0.583975mV 903075.756p 0.545934mV 904036.071p 0.577654mV 904039.185p 0.577654mV 904078.307p 0.639262mV 905001.249p 0.553905mV 905051.384p 0.600705mV 905063.962p 0.600498mV 905071.816p 0.60189mV 905085.821p 0.579426mV 905097.598p 0.582641mV 905109.386p 0.533759mV 905122.698p 0.565875mV 905134.677p 0.5704mV 905153.164p 0.6324mV 906009.056p 0.580703mV 906022.246p 0.503546mV 906051.412p 0.504601mV 906058.33p 0.477608mV 906067.057p 0.527892mV 906070.752p 0.499906mV 906088.854p 0.572378mV 906105.822p 0.563197mV 906115.055p 0.558262mV 906141.087p 0.520126mV 906161.131p 0.40282mV 906168.425p 0.424261mV 907014.62p 0.606351mV 907019.522p 0.580389mV 907063.109p 0.563359mV 907095.514p 0.552252mV 907096.786p 0.552252mV 907127.26p 0.465682mV 907152.957p 0.446458mV 907172.093p 0.338008mV 908003.376p 0.55146mV 908016.558p 0.525417mV 908071.938p 0.598796mV 908074.763p 0.598796mV 908086.788p 0.575281mV 909002.999p 0.553968mV 909032.612p 0.552162mV 909047.802p 0.579153mV 909061.398p 0.553612mV 909113.511p 0.48936mV 910015.529p 0.580897mV 910027.155p 0.531026mV 910054.627p 0.617976mV 910066.104p 0.652188mV 910089.59p 0.669384mV 911035.328p 0.470476mV 911083.83p 0.577441mV 911098.762p 0.644641mV 911104.1p 0.615504mV 911129.204p 0.633558mV 911174.09p 0.614736mV 911180.924p 0.619361mV 911183.521p 0.619361mV 911185.291p 0.59628mV 911244.552p 0.564197mV 911289.809p 0.478675mV 911326.544p 0.56005mV 911335.519p 0.514527mV 911351.318p 0.550128mV 911365.099p 0.5338mV 911401.835p 0.52791mV 911423.251p 0.586996mV 911428.885p 0.615101mV 911442.643p 0.543657mV 911523.35p 0.665839mV 911538.32p 0.748846mV 911547.485p 0.756348mV 912015.532p 0.572091mV 912040.411p 0.493421mV 912089.23p 0.503506mV 912091.05p 0.525558mV 912114.196p 0.559664mV 912118.047p 0.529017mV 913043.391p 0.618624mV 913044.471p 0.618624mV 914004.526p 0.552663mV 914005.409p 0.579998mV 914026.498p 0.638524mV 914035.765p 0.591652mV 914049.886p 0.54661mV 914070.307p 0.48586mV 914128.505p 0.353466mV 915003.615p 0.553388mV 915033.449p 0.659639mV 916012.766p 0.497108mV 916028.476p 0.523135mV 916044.766p 0.495128mV 916061.103p 0.434498mV 917013.827p 0.547352mV 917053.777p 0.498668mV 917096.964p 0.507343mV 917133.368p 0.50308mV 917133.699p 0.50308mV 918063.809p 0.669646mV 919024.222p 0.489524mV 919029.152p 0.461066mV 919054.202p 0.417943mV 920044.508p 0.42986mV 921028.605p 0.425815mV 922019.272p 0.629341mV 922030.584p 0.662362mV 922033.739p 0.662362mV 922039.645p 0.639628mV 923003.192p 0.553067mV 923064.526p 0.381878mV 924011.549p 0.495049mV 925120.799p 0.482106mV 926032.833p 0.542298mV 926042.282p 0.485381mV 926051.786p 0.532479mV 926061.511p 0.578432mV 926071.572p 0.572203mV 926096.348p 0.533379mV 926114.912p 0.500129mV 926120.684p 0.546104mV 926123.17p 0.546104mV 926128.98p 0.568727mV 926131.402p 0.591322mV 926161.974p 0.466973mV 926168.128p 0.436994mV 927007.385p 0.52362mV 927084.831p 0.47216mV 929004.004p 0.549849mV 929005.021p 0.524017mV 929041.83p 0.714222mV 929054.107p 0.668737mV 930024.271p 0.655445mV 930029.896p 0.682589mV 930032.48p 0.65776mV 930077.718p 0.614018mV 931010.415p 0.551143mV 931070.488p 0.542687mV 931094.727p 0.48058mV 931128.298p 0.530849mV 932000.86p 0.547444mV 932008.23p 0.521421mV 932023.873p 0.442595mV 932046.011p 0.460208mV 932066.768p 0.393074mV 933004.935p 0.553497mV 933015.131p 0.47044mV 933036.588p 0.459333mV 934041.599p 0.486116mV 934058.104p 0.399428mV 935014.303p 0.54878mV 935047.866p 0.522425mV 935048.57p 0.522425mV 935050.498p 0.494922mV 935062.405p 0.491875mV 935072.865p 0.540238mV 935075.642p 0.563989mV 936041.085p 0.608626mV 936053.521p 0.609731mV 936060.6p 0.559367mV 936081.682p 0.566259mV 936088.813p 0.542174mV 936114.622p 0.580755mV 936130.955p 0.489411mV 936147.191p 0.523602mV 936150.847p 0.49914mV 936184.289p 0.507402mV 936221.099p 0.569381mV 936223.367p 0.569381mV 936242.855p 0.576405mV 936243.282p 0.576405mV 936253.633p 0.579798mV 936308.924p 0.534587mV 936311.892p 0.511762mV 936326.596p 0.599372mV 936339.304p 0.605796mV 936355.549p 0.57107mV 936407.869p 0.566592mV 936408.492p 0.566592mV 936439.62p 0.541687mV 936462.44p 0.537853mV 936467.234p 0.567874mV 936467.948p 0.567874mV 937042.257p 0.496102mV 937069.313p 0.515162mV 937107.187p 0.437465mV 938108.992p 0.55916mV 938120.742p 0.568893mV 938120.833p 0.568893mV 938135.114p 0.527189mV 939003.828p 0.546105mV 939016.834p 0.523376mV 940002.034p 0.546584mV 940026.921p 0.686026mV 941006.328p 0.528694mV 941032.242p 0.559555mV 941051.829p 0.615196mV 941056.905p 0.642909mV 941082.117p 0.632703mV 942030.73p 0.649137mV 942035.037p 0.675622mV 942039.235p 0.675622mV 942041.965p 0.702716mV 942042.551p 0.702716mV 942062.067p 0.661409mV 942067.997p 0.639894mV 943020.036p 0.492137mV 943020.122p 0.492137mV 944009.929p 0.523792mV 944032.537p 0.437738mV 945011.919p 0.605147mV 945018.069p 0.632033mV 945022.688p 0.659254mV 945032.414p 0.610193mV 946021.322p 0.548835mV 946032.846p 0.601988mV 946048.098p 0.683291mV 946054.56p 0.65888mV 947025.191p 0.585401mV 947055.073p 0.501829mV 947083.905p 0.491701mV 947093.615p 0.54915mV 947099.28p 0.577543mV 947112.14p 0.610529mV 947113.624p 0.610529mV 947115.469p 0.586828mV 947134.243p 0.622537mV 947149.505p 0.609647mV 948045.635p 0.644098mV 948057.742p 0.652795mV 949002.757p 0.550794mV 949003.228p 0.550794mV 949035.979p 0.588148mV 949068.018p 0.657988mV 950021.797p 0.49867mV 950037.346p 0.522568mV 950037.552p 0.522568mV 950046.971p 0.466678mV 951006.082p 0.578484mV 951013.76p 0.552931mV 951018.159p 0.580212mV 951023.778p 0.554863mV 951047.017p 0.481444mV 951080.329p 0.451104mV 952028.962p 0.628385mV 952029.898p 0.628385mV 952074.208p 0.573413mV 952077.416p 0.551651mV 952090.146p 0.538743mV 952106.303p 0.524723mV 952128.037p 0.539537mV 952136.647p 0.49291mV 952137.311p 0.49291mV 952138.198p 0.49291mV 952152.725p 0.525876mV 952173.801p 0.531409mV 952198.97p 0.459441mV 952215.552p 0.458596mV 953038.71p 0.417639mV 953053.892p 0.489155mV 954005.042p 0.579731mV 954039.328p 0.483753mV 954095.887p 0.523684mV 954109.327p 0.464212mV 955012.16p 0.550224mV 955066.981p 0.456847mV 955069.814p 0.456847mV 956000.063p 0.549709mV 956042.478p 0.551641mV 956045.243p 0.526267mV 956073.004p 0.556624mV 956140.965p 0.454671mV 957000.959p 0.553442mV 957031.793p 0.663413mV 957033.423p 0.663413mV 958002.089p 0.55054mV 958038.735p 0.572826mV 958043.374p 0.598727mV 958059.335p 0.572263mV 958072.825p 0.652247mV 958076.675p 0.679612mV 958103.389p 0.563854mV 958116.915p 0.603106mV 959055.828p 0.571161mV 959079.641p 0.62582mV 959081.736p 0.600421mV 959081.758p 0.600421mV 959086.97p 0.575521mV 959090.795p 0.550958mV 959096.262p 0.579117mV 959128.956p 0.59444mV 960014.589p 0.548914mV 960030.987p 0.553256mV 960057.478p 0.480942mV 960097.106p 0.529427mV 960124.596p 0.604039mV 960128.352p 0.576937mV 960152.313p 0.604478mV 960155.99p 0.579924mV 960156.644p 0.579924mV 960188.459p 0.540642mV 960209.346p 0.549048mV 960224.108p 0.633362mV 960242.824p 0.646592mV 961012.304p 0.499135mV 961035.559p 0.623008mV 961036.532p 0.623008mV 961037.191p 0.623008mV 961063.695p 0.701656mV 962016.722p 0.576649mV 962018.762p 0.576649mV 962018.799p 0.576649mV 962026.908p 0.577143mV 962037.202p 0.630659mV 962045.068p 0.632867mV 962055.732p 0.584957mV 962063.543p 0.614057mV 962081.457p 0.576151mV 962087.261p 0.553979mV 962107.773p 0.518016mV 962130.432p 0.510645mV 962151.631p 0.470541mV 962165.549p 0.395021mV 963000.816p 0.552363mV 963010.761p 0.550537mV 963050.89p 0.438232mV 963051.482p 0.438232mV 964020.808p 0.605521mV 964026.981p 0.580671mV 964039.678p 0.584457mV 964071.166p 0.58156mV 964079.738p 0.560726mV 964081.775p 0.591776mV 965020.329p 0.601155mV 965029.232p 0.626618mV 965042.492p 0.599935mV 965047.215p 0.626675mV 965064.464p 0.603789mV 965069.467p 0.632067mV 965085.995p 0.592825mV 965091.911p 0.623285mV 965095.443p 0.653953mV 965097.103p 0.653953mV 966037.208p 0.521513mV 966073.252p 0.482157mV 967021.834p 0.504006mV 967076.179p 0.530757mV 967080.607p 0.504165mV 967086.308p 0.477453mV 967088.438p 0.477453mV 967093.911p 0.450459mV 967108.013p 0.471686mV 968028.091p 0.461269mV 968030.623p 0.432791mV 969013.619p 0.547967mV 969013.872p 0.547967mV 969034.568p 0.652319mV 969041.218p 0.654006mV 969062.121p 0.664246mV 970008.916p 0.526317mV 970009.322p 0.526317mV 970071.639p 0.606027mV 970076.683p 0.632494mV 970110.63p 0.61847mV 970132.249p 0.687036mV 971004.101p 0.548954mV 971017.215p 0.57323mV 971031.387p 0.545031mV 971034.581p 0.545031mV 971036.318p 0.571144mV 971044.921p 0.597225mV 971050.647p 0.597271mV 971066.212p 0.626584mV 971121.927p 0.641728mV 972006.549p 0.522905mV 972010.831p 0.496697mV 973012.699p 0.600246mV 973050.273p 0.666569mV 974023.493p 0.500403mV 974041.031p 0.496735mV 974079.006p 0.503192mV 975000.298p 0.552042mV 975048.406p 0.62346mV 975052.644p 0.596228mV 975054.371p 0.596228mV 975073.195p 0.64854mV 975104.248p 0.661042mV 976005.409p 0.579343mV 976020.137p 0.603334mV 976033.214p 0.603037mV 976043.531p 0.657074mV 976047.599p 0.684732mV 976053.942p 0.713008mV 977003.951p 0.550008mV 977044.489p 0.440486mV 977063.291p 0.323422mV 978002.257p 0.551857mV 978040.669p 0.444752mV 978040.993p 0.444752mV 978056.21p 0.410147mV 979030.822p 0.598911mV 979051.618p 0.651926mV 979066.338p 0.577603mV 979101.43p 0.629253mV 980050.936p 0.674292mV 980051.165p 0.674292mV 981012.396p 0.545697mV 981025.344p 0.515108mV 983015.914p 0.581609mV 983040.623p 0.511199mV 983078.606p 0.382464mV 984044.536p 0.539411mV 984045.179p 0.51109mV 984083.594p 0.519291mV 984100.124p 0.454427mV 985010.267p 0.545418mV 985062.841p 0.6481mV 985071.256p 0.703023mV 985085.102p 0.738326mV 986005.754p 0.577908mV 986047.208p 0.628421mV 986054.232p 0.603803mV 986068.873p 0.637684mV 986077.5p 0.697138mV 986078.769p 0.697138mV 987010.031p 0.547498mV 987069.584p 0.52851mV 987090.443p 0.452116mV 987093.747p 0.452116mV 987095.247p 0.477263mV 987130.36p 0.429978mV 988007.721p 0.521053mV 988028.169p 0.465549mV 988042.949p 0.433158mV 990023.98p 0.601529mV 990031.737p 0.603323mV 990043.152p 0.606126mV 990045.885p 0.581935mV 990049.757p 0.581935mV 990050.248p 0.610591mV 990087.345p 0.503158mV 990109.687p 0.568594mV 991009.637p 0.578042mV 991009.692p 0.578042mV 991034.492p 0.662021mV 992021.337p 0.603043mV 992023.825p 0.603043mV 992054.401p 0.563608mV 992066.393p 0.600843mV 992078.603p 0.661274mV 992084.091p 0.692012mV 993025.044p 0.517573mV 993051.027p 0.478745mV 994000.352p 0.549433mV 994000.615p 0.549433mV 994039.004p 0.46284mV 994039.82p 0.46284mV 995009.766p 0.521252mV 995039.127p 0.414751mV 995042.876p 0.386723mV 996011.955p 0.605649mV 996013.558p 0.605649mV 996014.142p 0.605649mV 996046.542p 0.541278mV 996078.036p 0.60824mV 996086.019p 0.665824mV 997027.631p 0.578199mV 997044.651p 0.501538mV 997061.228p 0.449519mV 998030.899p 0.595577mV 998039.64p 0.621548mV 998078.81p 0.691907mV 999008.147p 0.571106mV 999016.767p 0.516037mV 999028.789p 0.513443mV)
.ENDS conductors__anyBias-Lk_0_704



XVI1 28 285 conductors__anyBias-Lk_0_701
XREF1 B1 285 gnd newJTL__phaseReference
RR1  28 285 100

XVI2  37 385 conductors__anyBias-Lk_0_702
XREF2 B2 385 gnd newJTL__phaseReference
RR2  37 385 100

XVI3  64 485 conductors__anyBias-Lk_0_703
XREF3 B3 485 gnd newJTL__phaseReference
RR3  64 485 100

XVI4  73  585 conductors__anyBias-Lk_0_704
XREF4 B4 585 gnd newJTL__phaseReference
RR4 73  585  100






****TOP LEVEL CELL: aNewTestLibrary:testJTL{sch}


XJ1 1 junctionsBypassGround__gbj1p0
Xbias1 1 conductors__anyBias-Lk_0
XLL1 1 2 inductors__fixedInd1p5
XJ2 2 junctionsBypassGround__gbj1p0
Xbias2 2 conductors__anyBias-Lk_0
XLL2 2 3 inductors__fixedInd1p5
XJ3 3 junctionsBypassGround__gbj1p0
Xbias3 3 conductors__anyBias-Lk_0
XLL3 3 4 inductors__fixedInd1p5
XJ4 4 junctionsBypassGround__gbj1p0
Xbias4 4 conductors__anyBias-Lk_0
XLL4 4 5 inductors__fixedInd1p5
XJ5 5 junctionsBypassGround__gbj1p0
Xbias5 5 conductors__anyBias-Lk_0
XLL5 5 6 inductors__fixedInd1p5
XJ6 6 junctionsBypassGround__gbj1p0
Xbias6 6 conductors__anyBias-Lk_0
XLL6 6 7 inductors__fixedInd1p5
XJ7 7 junctionsBypassGround__gbj1p0
Xbias7 7 conductors__anyBias-Lk_0
XLL7 7 8 inductors__fixedInd1p5
XJ8 8 junctionsBypassGround__gbj1p0
Xbias8 8 conductors__anyBias-Lk_0
XLL8 8 9 inductors__fixedInd1p5
XJ9 9 junctionsBypassGround__gbj1p0
Xbias9 9 conductors__anyBias-Lk_0

XLL100 1 11 inductors__fixedInd1p5
XLL200 2 12 inductors__fixedInd1p5
XLL300 3 13 inductors__fixedInd1p5
XLL400 4 14 inductors__fixedInd1p5
XLL500 5 15 inductors__fixedInd1p5
XLL600 6 16 inductors__fixedInd1p5
XLL700 7 17 inductors__fixedInd1p5
XLL800 8 18 inductors__fixedInd1p5
XLL900 9 19 inductors__fixedInd1p5


XJ10 11 junctionsBypassGround__gbj1p0
Xbias10 11 conductors__anyBias-Lk_0
XLL10 11 12 inductors__fixedInd1p5
XJ11 12 junctionsBypassGround__gbj1p0
Xbias11 12 conductors__anyBias-Lk_0
XLL11 12 13 inductors__fixedInd1p5
XJ12 13 junctionsBypassGround__gbj1p0
Xbias12 13 conductors__anyBias-Lk_0
XLL12 13 14 inductors__fixedInd1p5
XJ13 14 junctionsBypassGround__gbj1p0
Xbias13 14 conductors__anyBias-Lk_0
XLL13 14 15 inductors__fixedInd1p5
XJ14 15 junctionsBypassGround__gbj1p0
Xbias14 15 conductors__anyBias-Lk_0
XLL14 15 16 inductors__fixedInd1p5
XJ15 16 junctionsBypassGround__gbj1p0
Xbias15 16 conductors__anyBias-Lk_0
XLL15 16 17 inductors__fixedInd1p5
XJ16 17 junctionsBypassGround__gbj1p0
Xbias16 17 conductors__anyBias-Lk_0
XLL16 17 18 inductors__fixedInd1p5
XJ17 18 junctionsBypassGround__gbj1p0
Xbias17 18 conductors__anyBias-Lk_0
XLL17 17 18 inductors__fixedInd1p5
XJ18 19 junctionsBypassGround__gbj1p0
Xbias18 19 conductors__anyBias-Lk_0

XLL110  11 21 inductors__fixedInd1p5
XLL210  12 22 inductors__fixedInd1p5
XLL310  13 23 inductors__fixedInd1p5
XLL410  14 24 inductors__fixedInd1p5
XLL510  15 25 inductors__fixedInd1p5
XLL610  16 26 inductors__fixedInd1p5
XLL710  17 27 inductors__fixedInd1p5
XLL810  18 28 inductors__fixedInd1p5
XLL910  19 29 inductors__fixedInd1p5

XJ19 21 junctionsBypassGround__gbj1p0
XLL19 21 22 inductors__fixedInd1p5
Xbias19 21 conductors__anyBias-Lk_0
XJ20 22 junctionsBypassGround__gbj1p0
Xbias20 22 conductors__anyBias-Lk_0
XLL20 22 23 inductors__fixedInd1p5
XJ21 23 junctionsBypassGround__gbj1p0
XLL21 23 24 inductors__fixedInd1p5
Xbias21 23 conductors__anyBias-Lk_0
XJ22 24 junctionsBypassGround__gbj1p0
Xbias22 24 conductors__anyBias-Lk_0
XLL22 24 25 inductors__fixedInd1p5
XJ23 25 junctionsBypassGround__gbj1p0
Xbias23 25 conductors__anyBias-Lk_0
XLL23 25 26 inductors__fixedInd1p5
XJ24 26 junctionsBypassGround__gbj1p0
Xbias24 26 conductors__anyBias-Lk_0
XLL24 26 27 inductors__fixedInd1p5
XJ25 27 junctionsBypassGround__gbj1p0
Xbias25 27 conductors__anyBias-Lk_0
XLL25 27 28 inductors__fixedInd1p5
XJ26 28 junctionsBypassGround__gbj1p0
Xbias26 28 conductors__anyBias-Lk_0
XLL26 28 29 inductors__fixedInd1p5
XJ27 29 junctionsBypassGround__gbj1p0
Xbias27 29 conductors__anyBias-Lk_0

XLL120   21 31 inductors__fixedInd1p5
XLL220   22 32 inductors__fixedInd1p5
XLL320   23 33 inductors__fixedInd1p5
XLL420   24 34 inductors__fixedInd1p5
XLL520   25 35 inductors__fixedInd1p5
XLL620   26 36 inductors__fixedInd1p5
XLL720   27 37 inductors__fixedInd1p5
XLL820   28 38 inductors__fixedInd1p5
XLL920   29 39 inductors__fixedInd1p5


XJ28 31 junctionsBypassGround__gbj1p0
XLL28 31 32 inductors__fixedInd1p5
Xbias28 31 conductors__anyBias-Lk_0
XJ29 32 junctionsBypassGround__gbj1p0
Xbias29 32 conductors__anyBias-Lk_0
XLL29 32 33 inductors__fixedInd1p5
XJ30 33 junctionsBypassGround__gbj1p0
XLL30 33 34 inductors__fixedInd1p5
Xbias30 33 conductors__anyBias-Lk_0
XJ31 34 junctionsBypassGround__gbj1p0
Xbias31 34 conductors__anyBias-Lk_0
XLL31 34 35 inductors__fixedInd1p5
XJ32 35 junctionsBypassGround__gbj1p0
Xbias32 35 conductors__anyBias-Lk_0
XLL32 35 36 inductors__fixedInd1p5
XJ33 36 junctionsBypassGround__gbj1p0
Xbias33 36 conductors__anyBias-Lk_0
XLL33 36 37 inductors__fixedInd1p5
XJ34 37 junctionsBypassGround__gbj1p0
Xbias34 37 conductors__anyBias-Lk_0
XLL34 37 38 inductors__fixedInd1p5
XJ35 38 junctionsBypassGround__gbj1p0
Xbias35 38 conductors__anyBias-Lk_0
XLL35 38 39 inductors__fixedInd1p5
XJ36 39 junctionsBypassGround__gbj1p0
Xbias36 39 conductors__anyBias-Lk_0


XLL130  31 41 inductors__fixedInd1p5
XLL230  32 42 inductors__fixedInd1p5
XLL330  33 43 inductors__fixedInd1p5
XLL430  34 44 inductors__fixedInd1p5
XLL530  35 45 inductors__fixedInd1p5
XLL630  36 46 inductors__fixedInd1p5
XLL730  37 47 inductors__fixedInd1p5
XLL830  38 48 inductors__fixedInd1p5
XLL930  39 49 inductors__fixedInd1p5



XJ37 41 junctionsBypassGround__gbj1p0
Xbias37 41 conductors__anyBias-Lk_0
XLL37 41 42 inductors__fixedInd1p5
XJ38 42 junctionsBypassGround__gbj1p0
Xbias38 42 conductors__anyBias-Lk_0
XLL38 42 43 inductors__fixedInd1p5
XJ39 43 junctionsBypassGround__gbj1p0
Xbias39 43 conductors__anyBias-Lk_0
XLL39 43 44 inductors__fixedInd1p5
XJ40 44 junctionsBypassGround__gbj1p0
Xbias40 44 conductors__anyBias-Lk_0
XLL40 44 45 inductors__fixedInd1p5
XJ41 45 junctionsBypassGround__gbj1p0
Xbias41 45 conductors__anyBias-Lk_0
XLL41 45 46 inductors__fixedInd1p5
XJ42 46 junctionsBypassGround__gbj1p0
Xbias42 46 conductors__anyBias-Lk_0
XLL42 46 47 inductors__fixedInd1p5
XJ43 47 junctionsBypassGround__gbj1p0
Xbias43 47 conductors__anyBias-Lk_0
XLL43 47 48 inductors__fixedInd1p5
XJ44 48 junctionsBypassGround__gbj1p0
Xbias44 48 conductors__anyBias-Lk_0
XLL44 48 49 inductors__fixedInd1p5
XJ45 49 junctionsBypassGround__gbj1p0
Xbias45 49 conductors__anyBias-Lk_0


XLL140  41 51 inductors__fixedInd1p5
XLL240  42 52 inductors__fixedInd1p5
XLL340  43 53 inductors__fixedInd1p5
XLL440  44 54 inductors__fixedInd1p5
XLL540  45 55 inductors__fixedInd1p5
XLL640  46 56 inductors__fixedInd1p5
XLL740  47 57 inductors__fixedInd1p5
XLL840  48 58 inductors__fixedInd1p5
XLL940  49 59 inductors__fixedInd1p5

XJ46 51 junctionsBypassGround__gbj1p0
Xbias46 51 conductors__anyBias-Lk_0
XLL46 51 52 inductors__fixedInd1p5
XJ47 52 junctionsBypassGround__gbj1p0
Xbias47 52 conductors__anyBias-Lk_0
XLL47 52 53 inductors__fixedInd1p5
XJ48 53 junctionsBypassGround__gbj1p0
Xbias48 53 conductors__anyBias-Lk_0
XLL48 53 54 inductors__fixedInd1p5
XJ49 54 junctionsBypassGround__gbj1p0
Xbias49 54 conductors__anyBias-Lk_0
XLL49 54 55 inductors__fixedInd1p5
XJ50 55 junctionsBypassGround__gbj1p0
Xbias50 55 conductors__anyBias-Lk_0
XLL50 55 56 inductors__fixedInd1p5
XJ51 56 junctionsBypassGround__gbj1p0
Xbias51 56 conductors__anyBias-Lk_0
XLL51 56 57 inductors__fixedInd1p5
XJ52 57 junctionsBypassGround__gbj1p0
Xbias52 57 conductors__anyBias-Lk_0
XLL52 57 58 inductors__fixedInd1p5
XJ53 58 junctionsBypassGround__gbj1p0
Xbias53 58 conductors__anyBias-Lk_0
XLL53 58 59 inductors__fixedInd1p5
XJ54 59 junctionsBypassGround__gbj1p0
Xbias54 59 conductors__anyBias-Lk_0

XLL150  51 61 inductors__fixedInd1p5
XLL250  52 62 inductors__fixedInd1p5
XLL350  53 63 inductors__fixedInd1p5
XLL450  54 64 inductors__fixedInd1p5
XLL550  55 65 inductors__fixedInd1p5
XLL650  56 66 inductors__fixedInd1p5
XLL750  57 67 inductors__fixedInd1p5
XLL850  58 68 inductors__fixedInd1p5
XLL950  59 69 inductors__fixedInd1p5

XJ55 61 junctionsBypassGround__gbj1p0
Xbias55 61 conductors__anyBias-Lk_0
XLL55 61 62 inductors__fixedInd1p5
XJ56 62 junctionsBypassGround__gbj1p0
Xbias56 62 conductors__anyBias-Lk_0
XLL56 62 63 inductors__fixedInd1p5
XJ57 63 junctionsBypassGround__gbj1p0
Xbias57 63 conductors__anyBias-Lk_0
XLL57 63 64 inductors__fixedInd1p5
XJ58 64 junctionsBypassGround__gbj1p0
Xbias58 64 conductors__anyBias-Lk_0
XLL58 64 65 inductors__fixedInd1p5
XJ59 65 junctionsBypassGround__gbj1p0
Xbias59 65 conductors__anyBias-Lk_0
XLL59 65 66 inductors__fixedInd1p5
XJ60 66 junctionsBypassGround__gbj1p0
Xbias60 66 conductors__anyBias-Lk_0
XLL60 66 67 inductors__fixedInd1p5
XJ61 67 junctionsBypassGround__gbj1p0
Xbias61 67 conductors__anyBias-Lk_0
XLL61 67 68 inductors__fixedInd1p5
XJ62 68 junctionsBypassGround__gbj1p0
Xbias62 68 conductors__anyBias-Lk_0
XLL62 68 69 inductors__fixedInd1p5
XJ63 69 junctionsBypassGround__gbj1p0
Xbias63 69 conductors__anyBias-Lk_0


XLL160  61 71 inductors__fixedInd1p5
XLL260  62 72 inductors__fixedInd1p5
XLL360  63 73 inductors__fixedInd1p5
XLL460  64 74 inductors__fixedInd1p5
XLL560  65 75 inductors__fixedInd1p5
XLL660  66 76 inductors__fixedInd1p5
XLL760  67 77 inductors__fixedInd1p5
XLL860  68 78 inductors__fixedInd1p5
XLL960  69 79 inductors__fixedInd1p5


XJ64 71 junctionsBypassGround__gbj1p0
Xbias64 71 conductors__anyBias-Lk_0
XLL64 71 72 inductors__fixedInd1p5
XJ65 72 junctionsBypassGround__gbj1p0
Xbias65 72 conductors__anyBias-Lk_0
XLL65 72 73 inductors__fixedInd1p5
XJ66 73 junctionsBypassGround__gbj1p0
Xbias66 73 conductors__anyBias-Lk_0
XLL66 73 74 inductors__fixedInd1p5
XJ67 74 junctionsBypassGround__gbj1p0
Xbias67 74 conductors__anyBias-Lk_0
XLL67 74 75 inductors__fixedInd1p5
XJ68 75 junctionsBypassGround__gbj1p0
Xbias68 75 conductors__anyBias-Lk_0
XLL68 75 76 inductors__fixedInd1p5
XJ69 76 junctionsBypassGround__gbj1p0
Xbias69 76 conductors__anyBias-Lk_0
XLL69 76 77 inductors__fixedInd1p5
XJ70 77 junctionsBypassGround__gbj1p0
Xbias70 77 conductors__anyBias-Lk_0
XLL70 77 78 inductors__fixedInd1p5
XJ71 78 junctionsBypassGround__gbj1p0
Xbias71 78 conductors__anyBias-Lk_0
XLL71 78 79 inductors__fixedInd1p5
XJ72 79 junctionsBypassGround__gbj1p0
Xbias72 79 conductors__anyBias-Lk_0


XLL170  71 81 inductors__fixedInd1p5
XLL270  72 82 inductors__fixedInd1p5
XLL370  73 83 inductors__fixedInd1p5
XLL470  74 84 inductors__fixedInd1p5
XLL570  75 85 inductors__fixedInd1p5
XLL670  76 86 inductors__fixedInd1p5
XLL770  77 87 inductors__fixedInd1p5
XLL870  78 88 inductors__fixedInd1p5
XLL970  79 89 inductors__fixedInd1p5


XJ73 81 junctionsBypassGround__gbj1p0
Xbias73 81 conductors__anyBias-Lk_0
XLL73 81 82 inductors__fixedInd1p5
XJ74 82 junctionsBypassGround__gbj1p0
Xbias74 82 conductors__anyBias-Lk_0
XLL74 82 83 inductors__fixedInd1p5
XJ75 83 junctionsBypassGround__gbj1p0
Xbias75 83 conductors__anyBias-Lk_0
XLL75 83 84 inductors__fixedInd1p5
XJ76 84 junctionsBypassGround__gbj1p0
Xbias76 84 conductors__anyBias-Lk_0
XLL76 84 85 inductors__fixedInd1p5
XJ77 85 junctionsBypassGround__gbj1p0
Xbias77 85 conductors__anyBias-Lk_0
XLL77 85 86 inductors__fixedInd1p5
XJ78 86 junctionsBypassGround__gbj1p0
Xbias78 86 conductors__anyBias-Lk_0
XLL78 86 87 inductors__fixedInd1p5
XJ79 87 junctionsBypassGround__gbj1p0
Xbias79 87 conductors__anyBias-Lk_0
XLL79 87 88 inductors__fixedInd1p5
XJ80 89 junctionsBypassGround__gbj1p0
Xbias80 89 conductors__anyBias-Lk_0
XLL80 89 90 inductors__fixedInd1p5
XJ81 91 junctionsBypassGround__gbj1p0
Xbias81 91 conductors__anyBias-Lk_0

.END
