*** SPICE deck for cell testJTLplain{sch} from library aNewTestLibrary
*** Created on Sat Jan 09, 2021 14:13:09
*** Last revised on Mon Aug 26, 2024 11:38:12
*** Written on Mon Aug 26, 2024 11:55:08 by Electric VLSI Design System, version 9.08e
*** Layout tech: josephson, foundry NONE
*** UC SPICE *** , MIN_RESIST 0.0, MIN_CAPAC 0.0FF
* Model cards copied from file: /Users/ivans/years/2020-2024/2024/2024-ivan/electric-2024/theBest1aug24/aTests/testJTLplain.txt
*** These are the print statement for testJTLplain
*** ies 26 August 2024
*** josim -o Aoutput.csv testJTLplain.cir 



.tran 0.1p 20p 0 0.1p


.print DEVI BJi|xJ40
.print DEVI BJi|xJ72
.print DEVI BJi|xJ33
.print DEVI BJi|xJ12
.print DEVI BJi|xJ73



* End of Model cards copied from file: /Users/ivans/years/2020-2024/2024/2024-ivan/electric-2024/theBest1jul24/aTests/testJTL.txt
.model jmitll jj(rtype=1, vg=.002V, cap=0.07pF, r0=160, rN=16, icrit=0.0001A)


.SUBCKT junctionsBypassGround__gbj1p0 D 
BJi D gnd jmitll area=1.25
RRi D gnd 5.36
.ENDS junctionsBypassGround__gbj1p0


*** SUBCIRCUIT inductors__fixedInd1p5 FROM CELL inductors:fixedInd3p0{sch}
.SUBCKT inductors__fixedInd1p5 A B
LLi A B 7.891E-12
.ENDS inductors__fixedInd1p5


*** SUBCIRCUIT conductors__anyBias-Lk_0 FROM CELL conductors:anyBias{sch}
.SUBCKT conductors__anyBias-Lk_0  D
RR1 NN D 29.42
VrampSppl@0 NN gnd pwl (0 0 1p 0.0026V)
.ENDS conductors__anyBias-Lk_0_707



****.SUBCKT conductors__anyBias-Lk_0 D
****RR1 NN D 8
****VrampSppl@0 NN gnd pwl (0 0 1p 3.86V)
***.ENDS conductors__anyBias-Lk_0

*** SUBCIRCUIT junctions__jb2p0 FROM CELL junctions:jb2p0{sch}
.SUBCKT junctions__jb2p0 D S
BJi S D jmitll area=2.5
RRi S D 2.68
.ENDS junctions__jb2p0

*** SUBCIRCUIT junctions__jb200p0 FROM CELL junctions:jb200p0{sch}
.SUBCKT junctions__jb200p0 D S
BJi S D jmitll area=250.0
RRi S D 0.0268
.ENDS junctions__jb200p0

*** SUBCIRCUIT conductors__anyBias-Lk_1_414 FROM CELL conductors:anyBias{sch}
.SUBCKT conductors__anyBias-Lk_1_414 D
RR1 NN D 14.71
VrampSppl@0 NN gnd pwl (0 0 1p 0.0026V)
.ENDS conductors__anyBias-Lk_1_414

*** SUBCIRCUIT conductors__bias1p4 FROM CELL conductors:bias1p4{sch}
.SUBCKT conductors__bias1p4 D
Xnormaliz@0 D conductors__anyBias-Lk_1_414
.ENDS conductors__bias1p4

*** SUBCIRCUIT conductors__anyBias-Lk_141_4 FROM CELL conductors:anyBias{sch}
.SUBCKT conductors__anyBias-Lk_141_4 D
RR1 NN D 0.147
VrampSppl@0 NN gnd pwl (0 0 1p 0.0026V)
.ENDS conductors__anyBias-Lk_141_4

*** SUBCIRCUIT conductors__bias1p4x100 FROM CELL conductors:bias1p4x100{sch}
.SUBCKT conductors__bias1p4x100 D
Xnormaliz@0 D conductors__anyBias-Lk_141_4
.ENDS conductors__bias1p4x100

*** SUBCIRCUIT newJTL__phaseReference FROM CELL newJTL:phaseReference{sch}
.SUBCKT newJTL__phaseReference B1 B2 gnd
XJ1 gnd B1 junctions__jb2p0
XJ2 gnd B2 junctions__jb200p0
LM1 net@4 B1 10e-16
LM2 net@3 B2 10e-16
Xbias1p4@0 net@4 conductors__bias1p4
Xbias1p4x@0 net@3 conductors__bias1p4x100
.ENDS newJTL__phaseReference







***Distorted3***
**.SUBCKT conductors__anyBias-Lk_0_701 bottom out
**VrampSppl@0 bottom out pwl (0 0 4.99p 0 5.0p 2mV 6p 2mV 6.1p 0 7.99p 0 8p 2mV 9p 2mV 9.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_701


**.SUBCKT conductors__anyBias-Lk_0_702 bottom out
**VrampSppl@0 bottom out pwl (0 0 10.9p 0 11p 2mV 12p 2mV 12.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_702

**.SUBCKT conductors__anyBias-Lk_0_703 bottom out
**VrampSppl@0 bottom out pwl (0 0 4.9p 0 5p 2mV 6p 2mV 6.1p 0 7.9p 0 8p 2mV 9p 2mV 9.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_703

**.SUBCKT conductors__anyBias-Lk_0_704  bottom out
**VrampSppl@0 bottom out pwl (0 0 10.9p 0 11p 2mV 12p 2mV 12.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_704

**.SUBCKT conductors__anyBias-Lk_0_705 bottom out
**VrampSppl@0 bottom out pwl (0 0 1.9p 0 2p 2mV 3p 2mV 3.1p 0 4.9p 0 5p 2mV 6p 2mV 6.1p 0 7.9p 0 8p 2mV 9p 2mV 9.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_705

***Distorted2***
**.SUBCKT conductors__anyBias-Lk_0_701 bottom out
**VrampSppl@0 bottom out pwl  (0 0 4.9p 0 5p 2mV 6p 2mV 6.1p 0 7.9p 0 8p 2mV 9p 2mV 9.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_701

**.SUBCKT conductors__anyBias-Lk_0_702 bottom out
**VrampSppl@0 bottom out pwl  (0 0 10.9p 0 11p 2mV 12p 2mV 12.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_702

**.SUBCKT conductors__anyBias-Lk_0_703 bottom out
**VrampSppl@0 bottom out pwl  (0 0 4.9p 0 5p 2mV 6p 2mV 6.1p 0 7.9p 0 8.0p 2mV 9p 2mV 9.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_703

**.SUBCKT conductors__anyBias-Lk_0_704 bottom out
**VrampSppl@0 bottom out pwl  (0 0 4.9p 0 5p 2mV 6p 2mV 6.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_704

**.SUBCKT conductors__anyBias-Lk_0_705 bottom out
**VrampSppl@0 bottom out pwl  (0 0 1.9p 0 2p 2mV 3p 2mV 3.1p 0 4.9p 0 5p 2mV 6p 2mV 6.1p 0 7.99p 0 8p 2mV 9p 2mV 9.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_705



**1**
**.SUBCKT conductors__anyBias-Lk_0_701 bottom out
**VrampSppl@0 bottom out pwl (0 0 7.9p 0 8p 2mV 9p 2mV 9.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_701


**.SUBCKT conductors__anyBias-Lk_0_702 bottom out
**VrampSppl@0 bottom out pwl (0 0 7.9p 0 8p 2mV 9p 2mV 9.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_702


**.SUBCKT conductors__anyBias-Lk_0_703 bottom out
**VrampSppl@0 bottom out pwl (0 0 7.9p 0 8p 2mV 9p 2mV 9.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_703

**.SUBCKT conductors__anyBias-Lk_0_704  bottom out
**VrampSppl@0 bottom out pwl  (0 0 7.9p 0 8p 2mV 9p 2mV 9.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_704

**.SUBCKT conductors__anyBias-Lk_0_705 bottom out
**VrampSppl@0 bottom out pwl (0 0 7.9p 0 8p 2mV 9p 2mV 9.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_705



***2***
**.SUBCKT conductors__anyBias-Lk_0_701 bottom out
**VrampSppl@0 bottom out pwl  (0 0 4.99p 0 5.0p 2mV 6p 2mV 6.1p 0 7.99p 0 8p 2mV 9p 2mV 9.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_701

**.SUBCKT conductors__anyBias-Lk_0_702 bottom out
**VrampSppl@0 bottom out pwl  (0 0 10.9p 0 11p 2mV 12p 2mV 12.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_702

**.SUBCKT conductors__anyBias-Lk_0_703 bottom out
**VrampSppl@0 bottom out pwl  (0 0 7.9p 0 8p 2mV 9p 2mV 10.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_703

**.SUBCKT conductors__anyBias-Lk_0_704 bottom out
**VrampSppl@0 bottom out pwl  (0 0 4.9p 0 5p 2mV 6p 2mV 7p 0p 15p 0)
**.ENDS conductors__anyBias-Lk_0_704

**.SUBCKT conductors__anyBias-Lk_0_705 bottom out
**VrampSppl@0 bottom out pwl  (0 0 1.9p 0 2p 2mV 3p 2mV 3.1p 0 4.9p 0 5.0p 2mV 6p 2mV 6.1p 0 7.99p 0 8p 2mV 9p 2mV 9.1p 0 10.9p 0 11p 2mV 12p 2mV 12.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_705

***3***
**.SUBCKT conductors__anyBias-Lk_0_701 bottom out
**VrampSppl@0 bottom out pwl (0 0 1.9p 0 2p 2mV 3p 2mV 3.1p 0 4.9p 0 5.0p 2mV 6p 2mV 6.1p 0 7.99p 0 8p 2mV 9p 2mV 9.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_701


**.SUBCKT conductors__anyBias-Lk_0_702 bottom out
**VrampSppl@0 bottom out pwl (0 0 10.9p 0 11p 2mV 12p 2mV 12.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_702

**.SUBCKT conductors__anyBias-Lk_0_703 bottom out
**VrampSppl@0 bottom out pwl (0 0 4.9p 0 5p 2mV 6p 2mV 6.1p 0 7.9p 0 8p 2mV 9p 2mV 9.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_703

**.SUBCKT conductors__anyBias-Lk_0_704  bottom out
**VrampSppl@0 bottom out pwl (0 0 10.9p 0 11p 2mV 12p 2mV 12.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_704

**.SUBCKT conductors__anyBias-Lk_0_705 bottom out
**VrampSppl@0 bottom out pwl (0 0 1.9p 0 2p 2mV 3p 2mV 3.1p 0 4.9p 0 5p 2mV 6p 2mV 6.1p 0 7.99p 0 8p 2mV 9p 2mV 9.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_705



***Distorted4***
**.SUBCKT conductors__anyBias-Lk_0_701 bottom out
**VrampSppl@0 bottom out pwl (0 0 4.9p 0 5p 2mV 6p 2mV 6.1p 0 7.9p 0 8p 2mV 9p 2mV 9.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_701


**.SUBCKT conductors__anyBias-Lk_0_702 bottom out
**VrampSppl@0 bottom out pwl (0 0 1.9p 0 2p 2mV 3p 2mV 3.1p 0 7.9p 0 8p 2mV 9p 2mV 9.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_702

**.SUBCKT conductors__anyBias-Lk_0_703 bottom out
**VrampSppl@0 bottom out pwl  (0 0 1.9p 0 2p 2mV 3p 2mV 3.1p 0 4.9p 0 5.0p 2mV 6p 2mV 6.1p 0 7.99p 0 8p 2mV 9p 2mV 9.1p 0 10.9p 0 11p 2mV 12p 2mV 12.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_703

**.SUBCKT conductors__anyBias-Lk_0_704  bottom out
**VrampSppl@0 bottom out pwl (0 0 7.9p 0 8p 2mV 9p 2mV 9.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_704

**.SUBCKT conductors__anyBias-Lk_0_705 bottom out
**VrampSppl@0 bottom out pwl (0 0 7.9p 0 8p 2mV 9p 2mV 9.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_705



***4***
**.SUBCKT conductors__anyBias-Lk_0_701 bottom out
**VrampSppl@0 bottom out pwl (0 0 1.9p 0 2p 2mV 3p 2mV 3.1p 0 7.9p 0 8p 2mV 9p 2mV 9.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_701


**.SUBCKT conductors__anyBias-Lk_0_702 bottom out
**VrampSppl@0 bottom out pwl (0 0 1.9p 0 2p 2mV 3p 2mV 3.1p 0 7.9p 0 8p 2mV 9p 2mV 9.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_702

**.SUBCKT conductors__anyBias-Lk_0_703 bottom out
**VrampSppl@0 bottom out pwl  (0 0 1.9p 0 2p 2mV 3p 2mV 3.1p 0 4.9p 0 5.0p 2mV 6p 2mV 6.1p 0 7.99p 0 8p 2mV 9p 2mV 9.1p 0 10.9p 0 11p 2mV 12p 2mV 12.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_703

**.SUBCKT conductors__anyBias-Lk_0_704  bottom out
**VrampSppl@0 bottom out pwl (0 0 7.9p 0 8p 2mV 9p 2mV 9.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_704

**.SUBCKT conductors__anyBias-Lk_0_705 bottom out
**VrampSppl@0 bottom out pwl (0 0 7.9p 0 8p 2mV 9p 2mV 9.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_705


**5**
**.SUBCKT conductors__anyBias-Lk_0_701 bottom out
**VrampSppl@0 bottom out pwl  (0 0 4.9p 0 5.0p 2mV 6p 2mV 6.1p 0 7.99p 0 8p 2mV 9p 2mV 9.1p 0 10.9p 0 11p 2mV 12p 2mV 12.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_701


**.SUBCKT conductors__anyBias-Lk_0_702 bottom out
**VrampSppl@0 bottom out pwl (0 0 4.9p 0 5p 2mV 6p 2mV 7p 0p 15p 0)
**.ENDS conductors__anyBias-Lk_0_702

**.SUBCKT conductors__anyBias-Lk_0_703 bottom out
**VrampSppl@0 bottom out pwl (0 0 4.9p 0 5.0p 2mV 6p 2mV 6.1p 0 7.99p 0 8p 2mV 9p 2mV 9.1p 0 10.9p 0 11p 2mV 12p 2mV 12.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_703

**.SUBCKT conductors__anyBias-Lk_0_704  bottom out
**VrampSppl@0 bottom out pwl  (0 0 10.9p 0 11p 2mV 12p 2mV 12.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_704

**.SUBCKT conductors__anyBias-Lk_0_705 bottom out
**VrampSppl@0 bottom out pwl (0 0 1.9p 0 2p 2mV 3p 2mV 3.1p 0 4.9p 0 5.0p 2mV 6p 2mV 6.1p 0 7.99p 0 8p 2mV 9p 2mV 9.1p 0 10.9p 0 11p 2mV 12p 2mV 12.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_705


**6**
**.SUBCKT conductors__anyBias-Lk_0_701 bottom out
**VrampSppl@0 bottom out pwl  (0 0 1.9p 0 2p 2mV 3p 2mV 3.1p 0 4.9p 0 5.0p 2mV 6p 2mV 6.1p 0 7.99p 0 8p 2mV 9p 2mV 9.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_701


**.SUBCKT conductors__anyBias-Lk_0_702 bottom out
**VrampSppl@0 bottom out pwl (0 0 1.9p 0 2p 2mV 3p 2mV 3.1p 0p 15p 0)
**.ENDS conductors__anyBias-Lk_0_702

**.SUBCKT conductors__anyBias-Lk_0_703 bottom out
**VrampSppl@0 bottom out pwl (0 0 1.9p 0 2p 2mV 3p 2mV 3.1p 0 4.9p 0 5.0p 2mV 6p 2mV 6.1p 0 7.99p 0 8p 2mV 9p 2mV 9.1p 0 10.9p 0 11p 2mV 12p 2mV 12.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_703

**.SUBCKT conductors__anyBias-Lk_0_704  bottom out
**VrampSppl@0 bottom out pwl  (0 0 1.9p 0 2p 2mV 3p 2mV 3.1p 0 10.9p 0  11p 2mV  12p 2mV 12.1 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_704

**.SUBCKT conductors__anyBias-Lk_0_705 bottom out
**VrampSppl@0 bottom out pwl (0 0 1.9p 0 2p 2mV 3p 2mV 3.1p 0 4.9p 0 5.0p 2mV 6p 2mV 6.1p 0 7.99p 0 8p 2mV 9p 2mV 9.1p 0 10.9p 0 11p 2mV 12p 2mV 12.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_705





**Distorted7**
**.SUBCKT conductors__anyBias-Lk_0_701 bottom out
**VrampSppl@0 bottom out pwl  (0 0 1.9p 0 2p 2mV 3p 2mV 3.1p 0 4.9p 0 5.0p 2mV 6p 2mV 6.1p 0 7.99p 0 8p 2mV 9p 2mV 9.1p 0 10.9p 0 11p 2mV 12p 2mV 12.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_701


**.SUBCKT conductors__anyBias-Lk_0_702 bottom out
**VrampSppl@0 bottom out pwl (0 0 10.9p 0 11p 2mV 12p 2mV 12.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_702

**.SUBCKT conductors__anyBias-Lk_0_703 bottom out
**VrampSppl@0 bottom out pwl (0 0 7.9p 0 8p 2mV 9p 2mV 9.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_703

**.SUBCKT conductors__anyBias-Lk_0_704  bottom out
**VrampSppl@0 bottom out pwl  (0 0 7.9p 0 8p 2mV 9p 2mV 9.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_704

**.SUBCKT conductors__anyBias-Lk_0_705 bottom out
**VrampSppl@0 bottom out pwl (0 0 4.9p 0 5p 2mV 6p 2mV 6.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_705




**7**
**.SUBCKT conductors__anyBias-Lk_0_701 bottom out
**VrampSppl@0 bottom out pwl  (0 0 1.9p 0 2p 2mV 3p 2mV 3.1p 0 4.9p 0 5.0p 2mV 6p 2mV 6.1p 0 7.99p 0 8p 2mV 9p 2mV 9.1p 0 10.9p 0 11p 2mV 12p 2mV 12.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_701


**.SUBCKT conductors__anyBias-Lk_0_702 bottom out
**VrampSppl@0 bottom out pwl (0 0 10.9p 0 11p 2mV 12p 2mV 12.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_702

**.SUBCKT conductors__anyBias-Lk_0_703 bottom out
**VrampSppl@0 bottom out pwl (0 0 7.9p 0 8p 2mV 9p 2mV 9.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_703

**.SUBCKT conductors__anyBias-Lk_0_704  bottom out
**VrampSppl@0 bottom out pwl  (0 0 7.9p 0 8p 2mV 9p 2mV 9.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_704

**.SUBCKT conductors__anyBias-Lk_0_705 bottom out
**VrampSppl@0 bottom out pwl (0 0 7.9p 0 8p 2mV 9p 2mV 9.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_705


**Distorted8**
**.SUBCKT conductors__anyBias-Lk_0_701 bottom out
**VrampSppl@0 bottom out pwl  (0 0 1.9p 0 2p 2mV 3p 2mV 3.1p 0 4.9p 0 5.0p 2mV 6p 2mV 6.1p 0 7.99p 0 8p 2mV 9p 2mV 9.1p 0 10.9p 0 11p 2mV 12p 2mV 12.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_701


**.SUBCKT conductors__anyBias-Lk_0_702 bottom out
**VrampSppl@0 bottom out pwl (0 0 1.9p 0 2p 2mV 3p 2mV 3.1p 0 10.9p 0  11p 2mV  12p 2mV 12.1 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_702

**.SUBCKT conductors__anyBias-Lk_0_703 bottom out
**VrampSppl@0 bottom out pwl (0 0 1.9p 0 2p 2mV 3p 2mV 3.1p 0 4.9p 0 5.0p 2mV 6p 2mV 6.1p 0 7.99p 0 8p 2mV 9p 2mV 9.1p 0 10.9p 0 11p 2mV 12p 2mV 12.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_703

**.SUBCKT conductors__anyBias-Lk_0_704  bottom out
**VrampSppl@0 bottom out pwl  (0 0 1.9p 0 2p 2mV 3p 2mV 3.1p 0 10.9p 0  11p 2mV  12p 2mV 12.1 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_704

**.SUBCKT conductors__anyBias-Lk_0_705 bottom out
**VrampSppl@0 bottom out pwl (0 0 10.9p 0 11p 2mV 12p 2mV 12.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_705


**8**
**.SUBCKT conductors__anyBias-Lk_0_701 bottom out
**VrampSppl@0 bottom out pwl  (0 0 1.9p 0 2p 2mV 3p 2mV 3.1p 0 4.9p 0 5.0p 2mV 6p 2mV 6.1p 0 7.99p 0 8p 2mV 9p 2mV 9.1p 0 10.9p 0 11p 2mV 12p 2mV 12.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_701


**.SUBCKT conductors__anyBias-Lk_0_702 bottom out
**VrampSppl@0 bottom out pwl (0 0 1.9p 0 2p 2mV 3p 2mV 3.1p 0 10.9p 0  11p 2mV  12p 2mV 12.1 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_702

**.SUBCKT conductors__anyBias-Lk_0_703 bottom out
**VrampSppl@0 bottom out pwl (0 0 1.9p 0 2p 2mV 3p 2mV 3.1p 0 4.9p 0 5.0p 2mV 6p 2mV 6.1p 0 7.99p 0 8p 2mV 9p 2mV 9.1p 0 10.9p 0 11p 2mV 12p 2mV 12.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_703

**.SUBCKT conductors__anyBias-Lk_0_704  bottom out
**VrampSppl@0 bottom out pwl  (0 0 1.9p 0 2p 2mV 3p 2mV 3.1p 0 10.9p 0  11p 2mV  12p 2mV 12.1 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_704

**.SUBCKT conductors__anyBias-Lk_0_705 bottom out
**VrampSppl@0 bottom out pwl (0 0 1.9p 0 2p 2mV 3p 2mV 3.1p 0 4.9p 0 5.0p 2mV 6p 2mV 6.1p 0 7.99p 0 8p 2mV 9p 2mV 9.1p 0 10.9p 0 11p 2mV 12p 2mV 12.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_705



**9**
**.SUBCKT conductors__anyBias-Lk_0_701 bottom out
**VrampSppl@0 bottom out pwl  (0 0 1.9p 0 2p 2mV 3p 2mV 3.1p 0 4.9p 0 5.0p 2mV 6p 2mV 6.1p 0 7.99p 0 8p 2mV 9p 2mV 9.1p 0 10.9p 0 11p 2mV 12p 2mV 12.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_701


**.SUBCKT conductors__anyBias-Lk_0_702 bottom out
**VrampSppl@0 bottom out pwl (0 0 1.9p 0 2p 2mV 3p 2mV 3.1p 0 10.9p 0  11p 2mV  12p 2mV 12.1 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_702

**.SUBCKT conductors__anyBias-Lk_0_703 bottom out
**VrampSppl@0 bottom out pwl (0 0 1.9p 0 2p 2mV 3p 2mV 3.1p 0 4.9p 0 5.0p 2mV 6p 2mV 6.1p 0 7.99p 0 8p 2mV 9p 2mV 9.1p 0 10.9p 0 11p 2mV 12p 2mV 12.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_703

**.SUBCKT conductors__anyBias-Lk_0_704  bottom out
**VrampSppl@0 bottom out pwl  (0 0 10.9p 0  11p 2mV  12p 2mV 12.1 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_704

**.SUBCKT conductors__anyBias-Lk_0_705  bottom out
**VrampSppl@0 bottom out pwl  (0 0 10.9p 0  11p 2mV  12p 2mV 12.1 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_705


**0**
**.SUBCKT conductors__anyBias-Lk_0_701 bottom out
**VrampSppl@0 bottom out pwl  (0 0 1.9p 0 2p 2mV 3p 2mV 3.1p 0 4.9p 0 5.0p 2mV 6p 2mV 6.1p 0 7.99p 0 8p 2mV 9p 2mV 9.1p 0 10.9p 0 11p 2mV 12p 2mV 12.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_701


**.SUBCKT conductors__anyBias-Lk_0_702 bottom out
**VrampSppl@0 bottom out pwl (0 0 1.9p 0 2p 2mV 3p 2mV 3.1p 0 10.9p 0  11p 2mV  12p 2mV 12.1 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_702

**.SUBCKT conductors__anyBias-Lk_0_703 bottom out
**VrampSppl@0 bottom out pwl (0 0 1.9p 0 2p 2mV 3p 2mV 3.1p 0 10.9p 0  11p 2mV  12p 2mV 12.1 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_703

**.SUBCKT conductors__anyBias-Lk_0_704 bottom out
**VrampSppl@0 bottom out pwl (0 0 1.9p 0 2p 2mV 3p 2mV 3.1p 0 10.9p 0  11p 2mV  12p 2mV 12.1 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_704

**.SUBCKT conductors__anyBias-Lk_0_705 bottom out
**VrampSppl@0 bottom out pwl  (0 0 1.9p 0 2p 2mV 3p 2mV 3.1p 0 4.9p 0 5.0p 2mV 6p 2mV 6.1p 0 7.99p 0 8p 2mV 9p 2mV 9.1p 0 10.9p 0 11p 2mV 12p 2mV 12.1p 0 15p 0)
**.ENDS conductors__anyBias-Lk_0_705

XVI 44 285 parity_check 
XREF B1 285 gnd newJTL__phaseReference
RR  44 285 100

**XVI1 44 285 conductors__anyBias-Lk_0_701
**XREF1 B1 285 gnd newJTL__phaseReference
**RR1  44 285 100

**XVI2  79 385 conductors__anyBias-Lk_0_702
**XREF2 B2 385 gnd newJTL__phaseReference
**RR2  79 385 100

**XVI3  36 485 conductors__anyBias-Lk_0_703
**XREF3 B3 485 gnd newJTL__phaseReference
**RR3  36 485 100

**XVI4  13  585 conductors__anyBias-Lk_0_704
**XREF4 B4 585 gnd newJTL__phaseReference
**RR4 13  585  100

**XVI5  81 685 conductors__anyBias-Lk_0_705
**XREF5 B5 685 gnd newJTL__phaseReference
**RR5  81 685 100




****TOP LEVEL CELL: aNewTestLibrary:testJTL{sch}


XJ1 1 junctionsBypassGround__gbj1p0
Xbias1 1 conductors__anyBias-Lk_0
XLL1 1 2 inductors__fixedInd1p5
XJ2 2 junctionsBypassGround__gbj1p0
Xbias2 2 conductors__anyBias-Lk_0
XLL2 2 3 inductors__fixedInd1p5
XJ3 3 junctionsBypassGround__gbj1p0
Xbias3 3 conductors__anyBias-Lk_0
XLL3 3 4 inductors__fixedInd1p5
XJ4 4 junctionsBypassGround__gbj1p0
Xbias4 4 conductors__anyBias-Lk_0
XLL4 4 5 inductors__fixedInd1p5
XJ5 5 junctionsBypassGround__gbj1p0
Xbias5 5 conductors__anyBias-Lk_0
XLL5 5 6 inductors__fixedInd1p5
XJ6 6 junctionsBypassGround__gbj1p0
Xbias6 6 conductors__anyBias-Lk_0
XLL6 6 7 inductors__fixedInd1p5
XJ7 7 junctionsBypassGround__gbj1p0
Xbias7 7 conductors__anyBias-Lk_0
XLL7 7 8 inductors__fixedInd1p5
XJ8 8 junctionsBypassGround__gbj1p0
Xbias8 8 conductors__anyBias-Lk_0
XLL8 8 9 inductors__fixedInd1p5
XJ9 9 junctionsBypassGround__gbj1p0
Xbias9 9 conductors__anyBias-Lk_0

XLL100 1 11 inductors__fixedInd1p5
XLL200 2 12 inductors__fixedInd1p5
XLL300 3 13 inductors__fixedInd1p5
XLL400 4 14 inductors__fixedInd1p5
XLL500 5 15 inductors__fixedInd1p5
XLL600 6 16 inductors__fixedInd1p5
XLL700 7 17 inductors__fixedInd1p5
XLL800 8 18 inductors__fixedInd1p5
XLL900 9 19 inductors__fixedInd1p5


XJ10 11 junctionsBypassGround__gbj1p0
Xbias10 11 conductors__anyBias-Lk_0
XLL10 11 12 inductors__fixedInd1p5
XJ11 12 junctionsBypassGround__gbj1p0
Xbias11 12 conductors__anyBias-Lk_0
XLL11 12 13 inductors__fixedInd1p5
XJ12 13 junctionsBypassGround__gbj1p0
Xbias12 13 conductors__anyBias-Lk_0
XLL12 13 14 inductors__fixedInd1p5
XJ13 14 junctionsBypassGround__gbj1p0
Xbias13 14 conductors__anyBias-Lk_0
XLL13 14 15 inductors__fixedInd1p5
XJ14 15 junctionsBypassGround__gbj1p0
Xbias14 15 conductors__anyBias-Lk_0
XLL14 15 16 inductors__fixedInd1p5
XJ15 16 junctionsBypassGround__gbj1p0
Xbias15 16 conductors__anyBias-Lk_0
XLL15 16 17 inductors__fixedInd1p5
XJ16 17 junctionsBypassGround__gbj1p0
Xbias16 17 conductors__anyBias-Lk_0
XLL16 17 18 inductors__fixedInd1p5
XJ17 18 junctionsBypassGround__gbj1p0
Xbias17 18 conductors__anyBias-Lk_0
XLL17 17 18 inductors__fixedInd1p5
XJ18 19 junctionsBypassGround__gbj1p0
Xbias18 19 conductors__anyBias-Lk_0

XLL110  11 21 inductors__fixedInd1p5
XLL210  12 22 inductors__fixedInd1p5
XLL310  13 23 inductors__fixedInd1p5
XLL410  14 24 inductors__fixedInd1p5
XLL510  15 25 inductors__fixedInd1p5
XLL610  16 26 inductors__fixedInd1p5
XLL710  17 27 inductors__fixedInd1p5
XLL810  18 28 inductors__fixedInd1p5
XLL910  19 29 inductors__fixedInd1p5

XJ19 21 junctionsBypassGround__gbj1p0
XLL19 21 22 inductors__fixedInd1p5
Xbias19 21 conductors__anyBias-Lk_0
XJ20 22 junctionsBypassGround__gbj1p0
Xbias20 22 conductors__anyBias-Lk_0
XLL20 22 23 inductors__fixedInd1p5
XJ21 23 junctionsBypassGround__gbj1p0
XLL21 23 24 inductors__fixedInd1p5
Xbias21 23 conductors__anyBias-Lk_0
XJ22 24 junctionsBypassGround__gbj1p0
Xbias22 24 conductors__anyBias-Lk_0
XLL22 24 25 inductors__fixedInd1p5
XJ23 25 junctionsBypassGround__gbj1p0
Xbias23 25 conductors__anyBias-Lk_0
XLL23 25 26 inductors__fixedInd1p5
XJ24 26 junctionsBypassGround__gbj1p0
Xbias24 26 conductors__anyBias-Lk_0
XLL24 26 27 inductors__fixedInd1p5
XJ25 27 junctionsBypassGround__gbj1p0
Xbias25 27 conductors__anyBias-Lk_0
XLL25 27 28 inductors__fixedInd1p5
XJ26 28 junctionsBypassGround__gbj1p0
Xbias26 28 conductors__anyBias-Lk_0
XLL26 28 29 inductors__fixedInd1p5
XJ27 29 junctionsBypassGround__gbj1p0
Xbias27 29 conductors__anyBias-Lk_0

XLL120   21 31 inductors__fixedInd1p5
XLL220   22 32 inductors__fixedInd1p5
XLL320   23 33 inductors__fixedInd1p5
XLL420   24 34 inductors__fixedInd1p5
XLL520   25 35 inductors__fixedInd1p5
XLL620   26 36 inductors__fixedInd1p5
XLL720   27 37 inductors__fixedInd1p5
XLL820   28 38 inductors__fixedInd1p5
XLL920   29 39 inductors__fixedInd1p5


XJ28 31 junctionsBypassGround__gbj1p0
XLL28 31 32 inductors__fixedInd1p5
Xbias28 31 conductors__anyBias-Lk_0
XJ29 32 junctionsBypassGround__gbj1p0
Xbias29 32 conductors__anyBias-Lk_0
XLL29 32 33 inductors__fixedInd1p5
XJ30 33 junctionsBypassGround__gbj1p0
XLL30 33 34 inductors__fixedInd1p5
Xbias30 33 conductors__anyBias-Lk_0
XJ31 34 junctionsBypassGround__gbj1p0
Xbias31 34 conductors__anyBias-Lk_0
XLL31 34 35 inductors__fixedInd1p5
XJ32 35 junctionsBypassGround__gbj1p0
Xbias32 35 conductors__anyBias-Lk_0
XLL32 35 36 inductors__fixedInd1p5
XJ33 36 junctionsBypassGround__gbj1p0
Xbias33 36 conductors__anyBias-Lk_0
XLL33 36 37 inductors__fixedInd1p5
XJ34 37 junctionsBypassGround__gbj1p0
Xbias34 37 conductors__anyBias-Lk_0
XLL34 37 38 inductors__fixedInd1p5
XJ35 38 junctionsBypassGround__gbj1p0
Xbias35 38 conductors__anyBias-Lk_0
XLL35 38 39 inductors__fixedInd1p5
XJ36 39 junctionsBypassGround__gbj1p0
Xbias36 39 conductors__anyBias-Lk_0


XLL130  31 41 inductors__fixedInd1p5
XLL230  32 42 inductors__fixedInd1p5
XLL330  33 43 inductors__fixedInd1p5
XLL430  34 44 inductors__fixedInd1p5
XLL530  35 45 inductors__fixedInd1p5
XLL630  36 46 inductors__fixedInd1p5
XLL730  37 47 inductors__fixedInd1p5
XLL830  38 48 inductors__fixedInd1p5
XLL930  39 49 inductors__fixedInd1p5



XJ37 41 junctionsBypassGround__gbj1p0
Xbias37 41 conductors__anyBias-Lk_0
XLL37 41 42 inductors__fixedInd1p5
XJ38 42 junctionsBypassGround__gbj1p0
Xbias38 42 conductors__anyBias-Lk_0
XLL38 42 43 inductors__fixedInd1p5
XJ39 43 junctionsBypassGround__gbj1p0
Xbias39 43 conductors__anyBias-Lk_0
XLL39 43 44 inductors__fixedInd1p5
XJ40 44 junctionsBypassGround__gbj1p0
Xbias40 44 conductors__anyBias-Lk_0
XLL40 44 45 inductors__fixedInd1p5
XJ41 45 junctionsBypassGround__gbj1p0
Xbias41 45 conductors__anyBias-Lk_0
XLL41 45 46 inductors__fixedInd1p5
XJ42 46 junctionsBypassGround__gbj1p0
Xbias42 46 conductors__anyBias-Lk_0
XLL42 46 47 inductors__fixedInd1p5
XJ43 47 junctionsBypassGround__gbj1p0
Xbias43 47 conductors__anyBias-Lk_0
XLL43 47 48 inductors__fixedInd1p5
XJ44 48 junctionsBypassGround__gbj1p0
Xbias44 48 conductors__anyBias-Lk_0
XLL44 48 49 inductors__fixedInd1p5
XJ45 49 junctionsBypassGround__gbj1p0
Xbias45 49 conductors__anyBias-Lk_0


XLL140  41 51 inductors__fixedInd1p5
XLL240  42 52 inductors__fixedInd1p5
XLL340  43 53 inductors__fixedInd1p5
XLL440  44 54 inductors__fixedInd1p5
XLL540  45 55 inductors__fixedInd1p5
XLL640  46 56 inductors__fixedInd1p5
XLL740  47 57 inductors__fixedInd1p5
XLL840  48 58 inductors__fixedInd1p5
XLL940  49 59 inductors__fixedInd1p5

XJ46 51 junctionsBypassGround__gbj1p0
Xbias46 51 conductors__anyBias-Lk_0
XLL46 51 52 inductors__fixedInd1p5
XJ47 52 junctionsBypassGround__gbj1p0
Xbias47 52 conductors__anyBias-Lk_0
XLL47 52 53 inductors__fixedInd1p5
XJ48 53 junctionsBypassGround__gbj1p0
Xbias48 53 conductors__anyBias-Lk_0
XLL48 53 54 inductors__fixedInd1p5
XJ49 54 junctionsBypassGround__gbj1p0
Xbias49 54 conductors__anyBias-Lk_0
XLL49 54 55 inductors__fixedInd1p5
XJ50 55 junctionsBypassGround__gbj1p0
Xbias50 55 conductors__anyBias-Lk_0
XLL50 55 56 inductors__fixedInd1p5
XJ51 56 junctionsBypassGround__gbj1p0
Xbias51 56 conductors__anyBias-Lk_0
XLL51 56 57 inductors__fixedInd1p5
XJ52 57 junctionsBypassGround__gbj1p0
Xbias52 57 conductors__anyBias-Lk_0
XLL52 57 58 inductors__fixedInd1p5
XJ53 58 junctionsBypassGround__gbj1p0
Xbias53 58 conductors__anyBias-Lk_0
XLL53 58 59 inductors__fixedInd1p5
XJ54 59 junctionsBypassGround__gbj1p0
Xbias54 59 conductors__anyBias-Lk_0

XLL150  51 61 inductors__fixedInd1p5
XLL250  52 62 inductors__fixedInd1p5
XLL350  53 63 inductors__fixedInd1p5
XLL450  54 64 inductors__fixedInd1p5
XLL550  55 65 inductors__fixedInd1p5
XLL650  56 66 inductors__fixedInd1p5
XLL750  57 67 inductors__fixedInd1p5
XLL850  58 68 inductors__fixedInd1p5
XLL950  59 69 inductors__fixedInd1p5

XJ55 61 junctionsBypassGround__gbj1p0
Xbias55 61 conductors__anyBias-Lk_0
XLL55 61 62 inductors__fixedInd1p5
XJ56 62 junctionsBypassGround__gbj1p0
Xbias56 62 conductors__anyBias-Lk_0
XLL56 62 63 inductors__fixedInd1p5
XJ57 63 junctionsBypassGround__gbj1p0
Xbias57 63 conductors__anyBias-Lk_0
XLL57 63 64 inductors__fixedInd1p5
XJ58 64 junctionsBypassGround__gbj1p0
Xbias58 64 conductors__anyBias-Lk_0
XLL58 64 65 inductors__fixedInd1p5
XJ59 65 junctionsBypassGround__gbj1p0
Xbias59 65 conductors__anyBias-Lk_0
XLL59 65 66 inductors__fixedInd1p5
XJ60 66 junctionsBypassGround__gbj1p0
Xbias60 66 conductors__anyBias-Lk_0
XLL60 66 67 inductors__fixedInd1p5
XJ61 67 junctionsBypassGround__gbj1p0
Xbias61 67 conductors__anyBias-Lk_0
XLL61 67 68 inductors__fixedInd1p5
XJ62 68 junctionsBypassGround__gbj1p0
Xbias62 68 conductors__anyBias-Lk_0
XLL62 68 69 inductors__fixedInd1p5
XJ63 69 junctionsBypassGround__gbj1p0
Xbias63 69 conductors__anyBias-Lk_0


XLL160  61 71 inductors__fixedInd1p5
XLL260  62 72 inductors__fixedInd1p5
XLL360  63 73 inductors__fixedInd1p5
XLL460  64 74 inductors__fixedInd1p5
XLL560  65 75 inductors__fixedInd1p5
XLL660  66 76 inductors__fixedInd1p5
XLL760  67 77 inductors__fixedInd1p5
XLL860  68 78 inductors__fixedInd1p5
XLL960  69 79 inductors__fixedInd1p5


XJ64 71 junctionsBypassGround__gbj1p0
Xbias64 71 conductors__anyBias-Lk_0
XLL64 71 72 inductors__fixedInd1p5
XJ65 72 junctionsBypassGround__gbj1p0
Xbias65 72 conductors__anyBias-Lk_0
XLL65 72 73 inductors__fixedInd1p5
XJ66 73 junctionsBypassGround__gbj1p0
Xbias66 73 conductors__anyBias-Lk_0
XLL66 73 74 inductors__fixedInd1p5
XJ67 74 junctionsBypassGround__gbj1p0
Xbias67 74 conductors__anyBias-Lk_0
XLL67 74 75 inductors__fixedInd1p5
XJ68 75 junctionsBypassGround__gbj1p0
Xbias68 75 conductors__anyBias-Lk_0
XLL68 75 76 inductors__fixedInd1p5
XJ69 76 junctionsBypassGround__gbj1p0
Xbias69 76 conductors__anyBias-Lk_0
XLL69 76 77 inductors__fixedInd1p5
XJ70 77 junctionsBypassGround__gbj1p0
Xbias70 77 conductors__anyBias-Lk_0
XLL70 77 78 inductors__fixedInd1p5
XJ71 78 junctionsBypassGround__gbj1p0
Xbias71 78 conductors__anyBias-Lk_0
XLL71 78 79 inductors__fixedInd1p5
XJ72 79 junctionsBypassGround__gbj1p0
Xbias72 79 conductors__anyBias-Lk_0


XLL170  71 81 inductors__fixedInd1p5
XLL270  72 82 inductors__fixedInd1p5
XLL370  73 83 inductors__fixedInd1p5
XLL470  74 84 inductors__fixedInd1p5
XLL570  75 85 inductors__fixedInd1p5
XLL670  76 86 inductors__fixedInd1p5
XLL770  77 87 inductors__fixedInd1p5
XLL870  78 88 inductors__fixedInd1p5
XLL970  79 89 inductors__fixedInd1p5


XJ73 81 junctionsBypassGround__gbj1p0
Xbias73 81 conductors__anyBias-Lk_0
XLL73 81 82 inductors__fixedInd1p5
XJ74 82 junctionsBypassGround__gbj1p0
Xbias74 82 conductors__anyBias-Lk_0
XLL74 82 83 inductors__fixedInd1p5
XJ75 83 junctionsBypassGround__gbj1p0
Xbias75 83 conductors__anyBias-Lk_0
XLL75 83 84 inductors__fixedInd1p5
XJ76 84 junctionsBypassGround__gbj1p0
Xbias76 84 conductors__anyBias-Lk_0
XLL76 84 85 inductors__fixedInd1p5
XJ77 85 junctionsBypassGround__gbj1p0
Xbias77 85 conductors__anyBias-Lk_0
XLL77 85 86 inductors__fixedInd1p5
XJ78 86 junctionsBypassGround__gbj1p0
Xbias78 86 conductors__anyBias-Lk_0
XLL78 86 87 inductors__fixedInd1p5
XJ79 87 junctionsBypassGround__gbj1p0
Xbias79 87 conductors__anyBias-Lk_0
XLL79 87 88 inductors__fixedInd1p5
XJ80 89 junctionsBypassGround__gbj1p0
Xbias80 89 conductors__anyBias-Lk_0
XLL80 89 90 inductors__fixedInd1p5
XJ81 91 junctionsBypassGround__gbj1p0
Xbias81 91 conductors__anyBias-Lk_0

.END
